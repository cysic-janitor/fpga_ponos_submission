// --------------------------------------------------------------------------------
`timescale 1 ps / 1 ps

(* ORIG_REF_NAME = "shiftreg" *) 
module ponos_shiftreg
   (\DELAY_BLOCK[3].shift_array_reg[4] ,
    clk,
    prsi_red_scalar_i);
  output \DELAY_BLOCK[3].shift_array_reg[4] ;
  input clk;
  input [0:0]prsi_red_scalar_i;

  wire \<const0> ;
  wire \<const1> ;
  wire \DELAY_BLOCK[3].shift_array_reg[4] ;
  wire calc_add_sub_i;
  wire clk;
  wire [0:0]prsi_red_scalar_i;

  (* srl_bus_name = "\\i_shiftreg_calc_add_sub/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_add_sub/DELAY_BLOCK[3].shift_array_reg[4][0]_srl4 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][0]_srl4 
       (.A0(\<const1> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(calc_add_sub_i),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4] ));
  LUT1 #(
    .INIT(2'h1)) 
    \DELAY_BLOCK[3].shift_array_reg[4][0]_srl4_i_1 
       (.I0(prsi_red_scalar_i),
        .O(calc_add_sub_i));
  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
endmodule

(* ORIG_REF_NAME = "shiftreg" *) 
module ponos_shiftreg_0
   (calc_is_dummy_dld,
    clk,
    prsi_index_i);
  output calc_is_dummy_dld;
  input clk;
  input [2:0]prsi_index_i;

  wire \<const0> ;
  wire \<const1> ;
  wire \DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ;
  wire calc_is_dummy;
  wire calc_is_dummy_dld;
  wire clk;
  wire [2:0]prsi_index_i;

  (* srl_bus_name = "\\i_shiftreg_calc_is_dummy/DELAY_BLOCK[2].shift_array_reg[3] " *) 
  (* srl_name = "\\i_shiftreg_calc_is_dummy/DELAY_BLOCK[2].shift_array_reg[3][0]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[2].shift_array_reg[3][0]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(calc_is_dummy),
        .Q(\DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_i_1 
       (.I0(prsi_index_i[0]),
        .I1(prsi_index_i[1]),
        .I2(prsi_index_i[2]),
        .O(calc_is_dummy));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[3].shift_array_reg[4][0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ),
        .Q(calc_is_dummy_dld),
        .R(\<const0> ));
  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
endmodule

(* ORIG_REF_NAME = "shiftreg" *) 
module ponos_shiftreg_1
   (calc_is_zero_dld,
    \DELAY_BLOCK[3].shift_array_reg[4][0]_0 ,
    \DELAY_BLOCK[3].shift_array_reg[4][0]_1 ,
    \DELAY_BLOCK[3].shift_array_reg[4][0]_2 ,
    \DELAY_BLOCK[3].shift_array_reg[4][0]_3 ,
    \DELAY_BLOCK[3].shift_array_reg[4][0]_4 ,
    acc_valid_o0,
    calc_is_zero,
    clk,
    calc_is_dummy_dld,
    \accept_flags_o_reg[6] ,
    processing_first_accept_flag,
    Q,
    accept_flags_o,
    \accept_flags_o_reg[4] ,
    \accept_flags_o_reg[3] ,
    \accept_flags_o_reg[1] ,
    douta);
  output calc_is_zero_dld;
  output \DELAY_BLOCK[3].shift_array_reg[4][0]_0 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][0]_1 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][0]_2 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][0]_3 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][0]_4 ;
  output acc_valid_o0;
  input calc_is_zero;
  input clk;
  input calc_is_dummy_dld;
  input \accept_flags_o_reg[6] ;
  input processing_first_accept_flag;
  input [0:0]Q;
  input [3:0]accept_flags_o;
  input \accept_flags_o_reg[4] ;
  input \accept_flags_o_reg[3] ;
  input \accept_flags_o_reg[1] ;
  input [0:0]douta;

  wire \<const0> ;
  wire \<const1> ;
  wire \DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][0]_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][0]_1 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][0]_2 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][0]_3 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][0]_4 ;
  wire [0:0]Q;
  wire acc_valid_o0;
  wire [3:0]accept_flags_o;
  wire \accept_flags_o_reg[1] ;
  wire \accept_flags_o_reg[3] ;
  wire \accept_flags_o_reg[4] ;
  wire \accept_flags_o_reg[6] ;
  wire calc_is_dummy_dld;
  wire calc_is_zero;
  wire calc_is_zero_dld;
  wire clk;
  wire [0:0]douta;
  wire processing_first_accept_flag;

  (* srl_bus_name = "\\i_shiftreg_calc_is_zero/DELAY_BLOCK[2].shift_array_reg[3] " *) 
  (* srl_name = "\\i_shiftreg_calc_is_zero/DELAY_BLOCK[2].shift_array_reg[3][0]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[2].shift_array_reg[3][0]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(calc_is_zero),
        .Q(\DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[3].shift_array_reg[4][0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ),
        .Q(calc_is_zero_dld),
        .R(\<const0> ));
  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    acc_valid_o_i_1
       (.I0(Q),
        .I1(calc_is_zero_dld),
        .I2(douta),
        .I3(calc_is_dummy_dld),
        .O(acc_valid_o0));
  LUT6 #(
    .INIT(64'hFEFEFFFFFECE0000)) 
    \accept_flags_o[1]_i_1 
       (.I0(\DELAY_BLOCK[3].shift_array_reg[4][0]_1 ),
        .I1(calc_is_dummy_dld),
        .I2(\accept_flags_o_reg[1] ),
        .I3(processing_first_accept_flag),
        .I4(Q),
        .I5(accept_flags_o[0]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][0]_4 ));
  LUT6 #(
    .INIT(64'hFEFEFFFFFECE0000)) 
    \accept_flags_o[3]_i_1 
       (.I0(\DELAY_BLOCK[3].shift_array_reg[4][0]_1 ),
        .I1(calc_is_dummy_dld),
        .I2(\accept_flags_o_reg[3] ),
        .I3(processing_first_accept_flag),
        .I4(Q),
        .I5(accept_flags_o[1]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][0]_3 ));
  LUT6 #(
    .INIT(64'hFEFEFFFFFECE0000)) 
    \accept_flags_o[4]_i_1 
       (.I0(\DELAY_BLOCK[3].shift_array_reg[4][0]_1 ),
        .I1(calc_is_dummy_dld),
        .I2(\accept_flags_o_reg[4] ),
        .I3(processing_first_accept_flag),
        .I4(Q),
        .I5(accept_flags_o[2]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][0]_2 ));
  LUT6 #(
    .INIT(64'hFEFEFFFFFECE0000)) 
    \accept_flags_o[6]_i_1 
       (.I0(\DELAY_BLOCK[3].shift_array_reg[4][0]_1 ),
        .I1(calc_is_dummy_dld),
        .I2(\accept_flags_o_reg[6] ),
        .I3(processing_first_accept_flag),
        .I4(Q),
        .I5(accept_flags_o[3]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][0]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \accept_flags_o[6]_i_2 
       (.I0(calc_is_zero_dld),
        .I1(douta),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][0]_1 ));
endmodule

(* ORIG_REF_NAME = "shiftreg" *) 
module ponos_shiftreg__parameterized0
   (D,
    calc_is_zero,
    .prsi_red_scalar_i_4_sp_1(prsi_red_scalar_i_4_sn_1),
    data0,
    clk,
    prsi_red_scalar_i);
  output [11:0]D;
  output calc_is_zero;
  output [11:0]data0;
  input clk;
  input [12:0]prsi_red_scalar_i;
  output prsi_red_scalar_i_4_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [11:0]D;
  wire GND_2;
  wire calc_is_zero;
  wire clk;
  wire [11:0]data0;
  wire [12:0]prsi_red_scalar_i;
  wire prsi_red_scalar_i_4_sn_1;
  wire \shift_array[1][11]_i_10_n_0 ;
  wire \shift_array[1][11]_i_11_n_0 ;
  wire \shift_array[1][11]_i_12_n_0 ;
  wire \shift_array[1][11]_i_4_n_0 ;
  wire \shift_array[1][11]_i_5_n_0 ;
  wire \shift_array[1][11]_i_6_n_0 ;
  wire \shift_array[1][11]_i_7_n_0 ;
  wire \shift_array[1][11]_i_8_n_0 ;
  wire \shift_array[1][11]_i_9_n_0 ;
  wire \shift_array[1][7]_i_10_n_0 ;
  wire \shift_array[1][7]_i_11_n_0 ;
  wire \shift_array[1][7]_i_12_n_0 ;
  wire \shift_array[1][7]_i_13_n_0 ;
  wire \shift_array[1][7]_i_14_n_0 ;
  wire \shift_array[1][7]_i_15_n_0 ;
  wire \shift_array[1][7]_i_16_n_0 ;
  wire \shift_array[1][7]_i_17_n_0 ;
  wire \shift_array[1][7]_i_2_n_0 ;
  wire \shift_array[1][7]_i_3_n_0 ;
  wire \shift_array[1][7]_i_4_n_0 ;
  wire \shift_array[1][7]_i_5_n_0 ;
  wire \shift_array[1][7]_i_6_n_0 ;
  wire \shift_array[1][7]_i_7_n_0 ;
  wire \shift_array[1][7]_i_8_n_0 ;
  wire \shift_array[1][7]_i_9_n_0 ;
  wire \shift_array_reg[1][11]_i_2_n_5 ;
  wire \shift_array_reg[1][11]_i_2_n_6 ;
  wire \shift_array_reg[1][11]_i_2_n_7 ;
  wire \shift_array_reg[1][7]_i_1_n_0 ;
  wire \shift_array_reg[1][7]_i_1_n_1 ;
  wire \shift_array_reg[1][7]_i_1_n_2 ;
  wire \shift_array_reg[1][7]_i_1_n_3 ;
  wire \shift_array_reg[1][7]_i_1_n_4 ;
  wire \shift_array_reg[1][7]_i_1_n_5 ;
  wire \shift_array_reg[1][7]_i_1_n_6 ;
  wire \shift_array_reg[1][7]_i_1_n_7 ;
  wire \shift_array_reg_n_0_[1][0] ;
  wire \shift_array_reg_n_0_[1][10] ;
  wire \shift_array_reg_n_0_[1][11] ;
  wire \shift_array_reg_n_0_[1][1] ;
  wire \shift_array_reg_n_0_[1][2] ;
  wire \shift_array_reg_n_0_[1][3] ;
  wire \shift_array_reg_n_0_[1][4] ;
  wire \shift_array_reg_n_0_[1][5] ;
  wire \shift_array_reg_n_0_[1][6] ;
  wire \shift_array_reg_n_0_[1][7] ;
  wire \shift_array_reg_n_0_[1][8] ;
  wire \shift_array_reg_n_0_[1][9] ;

  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][0]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][0]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][0] ),
        .Q(D[0]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][10]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][10]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][10] ),
        .Q(D[10]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][11]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][11]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][11] ),
        .Q(D[11]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][1]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1] ),
        .Q(D[1]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][2]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][2]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][2] ),
        .Q(D[2]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][3]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][3]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][3] ),
        .Q(D[3]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][4]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][4]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][4] ),
        .Q(D[4]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][5]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][5]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][5] ),
        .Q(D[5]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][6]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][6]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][6] ),
        .Q(D[6]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][7]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][7]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][7] ),
        .Q(D[7]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][8]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][8]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][8] ),
        .Q(D[8]));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_addr/DELAY_BLOCK[3].shift_array_reg[4][9]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][9]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][9] ),
        .Q(D[9]));
  GND GND
       (.G(\<const0> ));
  GND GND_1
       (.G(GND_2));
  VCC VCC
       (.P(\<const1> ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][11]_i_1 
       (.I0(prsi_red_scalar_i_4_sn_1),
        .O(calc_is_zero));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][11]_i_10 
       (.I0(prsi_red_scalar_i[8]),
        .O(\shift_array[1][11]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \shift_array[1][11]_i_11 
       (.I0(prsi_red_scalar_i[8]),
        .I1(prsi_red_scalar_i[7]),
        .I2(prsi_red_scalar_i[10]),
        .I3(prsi_red_scalar_i[9]),
        .O(\shift_array[1][11]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \shift_array[1][11]_i_12 
       (.I0(prsi_red_scalar_i[0]),
        .I1(prsi_red_scalar_i[11]),
        .I2(prsi_red_scalar_i[12]),
        .I3(prsi_red_scalar_i[2]),
        .I4(prsi_red_scalar_i[1]),
        .O(\shift_array[1][11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \shift_array[1][11]_i_3 
       (.I0(\shift_array[1][11]_i_11_n_0 ),
        .I1(prsi_red_scalar_i[4]),
        .I2(prsi_red_scalar_i[3]),
        .I3(prsi_red_scalar_i[6]),
        .I4(prsi_red_scalar_i[5]),
        .I5(\shift_array[1][11]_i_12_n_0 ),
        .O(prsi_red_scalar_i_4_sn_1));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][11]_i_4 
       (.I0(prsi_red_scalar_i[10]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][11]_i_5 
       (.I0(prsi_red_scalar_i[9]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][11]_i_6 
       (.I0(prsi_red_scalar_i[8]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][11]_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][11]_i_7 
       (.I0(prsi_red_scalar_i[11]),
        .O(\shift_array[1][11]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][11]_i_8 
       (.I0(prsi_red_scalar_i[10]),
        .O(\shift_array[1][11]_i_8_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][11]_i_9 
       (.I0(prsi_red_scalar_i[9]),
        .O(\shift_array[1][11]_i_9_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][7]_i_10 
       (.I0(prsi_red_scalar_i[7]),
        .O(\shift_array[1][7]_i_10_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][7]_i_11 
       (.I0(prsi_red_scalar_i[6]),
        .O(\shift_array[1][7]_i_11_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][7]_i_12 
       (.I0(prsi_red_scalar_i[5]),
        .O(\shift_array[1][7]_i_12_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][7]_i_13 
       (.I0(prsi_red_scalar_i[4]),
        .O(\shift_array[1][7]_i_13_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][7]_i_14 
       (.I0(prsi_red_scalar_i[3]),
        .O(\shift_array[1][7]_i_14_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][7]_i_15 
       (.I0(prsi_red_scalar_i[2]),
        .O(\shift_array[1][7]_i_15_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][7]_i_16 
       (.I0(prsi_red_scalar_i[1]),
        .O(\shift_array[1][7]_i_16_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \shift_array[1][7]_i_17 
       (.I0(prsi_red_scalar_i[0]),
        .O(\shift_array[1][7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][7]_i_2 
       (.I0(prsi_red_scalar_i[7]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][7]_i_3 
       (.I0(prsi_red_scalar_i[6]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][7]_i_4 
       (.I0(prsi_red_scalar_i[5]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][7]_i_5 
       (.I0(prsi_red_scalar_i[4]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][7]_i_6 
       (.I0(prsi_red_scalar_i[3]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][7]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][7]_i_7 
       (.I0(prsi_red_scalar_i[2]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][7]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][7]_i_8 
       (.I0(prsi_red_scalar_i[1]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \shift_array[1][7]_i_9 
       (.I0(prsi_red_scalar_i[0]),
        .I1(prsi_red_scalar_i[12]),
        .O(\shift_array[1][7]_i_9_n_0 ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[0]),
        .Q(\shift_array_reg_n_0_[1][0] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[10]),
        .Q(\shift_array_reg_n_0_[1][10] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[11]),
        .Q(\shift_array_reg_n_0_[1][11] ),
        .R(calc_is_zero));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \shift_array_reg[1][11]_i_2 
       (.CI(\shift_array_reg[1][7]_i_1_n_0 ),
        .CI_TOP(GND_2),
        .CO({\shift_array_reg[1][11]_i_2_n_5 ,\shift_array_reg[1][11]_i_2_n_6 ,\shift_array_reg[1][11]_i_2_n_7 }),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\shift_array[1][11]_i_4_n_0 ,\shift_array[1][11]_i_5_n_0 ,\shift_array[1][11]_i_6_n_0 }),
        .O(data0[11:8]),
        .S({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\shift_array[1][11]_i_7_n_0 ,\shift_array[1][11]_i_8_n_0 ,\shift_array[1][11]_i_9_n_0 ,\shift_array[1][11]_i_10_n_0 }));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[1]),
        .Q(\shift_array_reg_n_0_[1][1] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[2]),
        .Q(\shift_array_reg_n_0_[1][2] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[3]),
        .Q(\shift_array_reg_n_0_[1][3] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[4]),
        .Q(\shift_array_reg_n_0_[1][4] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[5]),
        .Q(\shift_array_reg_n_0_[1][5] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[6]),
        .Q(\shift_array_reg_n_0_[1][6] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[7]),
        .Q(\shift_array_reg_n_0_[1][7] ),
        .R(calc_is_zero));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY8 #(
    .CARRY_TYPE("SINGLE_CY8")) 
    \shift_array_reg[1][7]_i_1 
       (.CI(\<const0> ),
        .CI_TOP(GND_2),
        .CO({\shift_array_reg[1][7]_i_1_n_0 ,\shift_array_reg[1][7]_i_1_n_1 ,\shift_array_reg[1][7]_i_1_n_2 ,\shift_array_reg[1][7]_i_1_n_3 ,\shift_array_reg[1][7]_i_1_n_4 ,\shift_array_reg[1][7]_i_1_n_5 ,\shift_array_reg[1][7]_i_1_n_6 ,\shift_array_reg[1][7]_i_1_n_7 }),
        .DI({\shift_array[1][7]_i_2_n_0 ,\shift_array[1][7]_i_3_n_0 ,\shift_array[1][7]_i_4_n_0 ,\shift_array[1][7]_i_5_n_0 ,\shift_array[1][7]_i_6_n_0 ,\shift_array[1][7]_i_7_n_0 ,\shift_array[1][7]_i_8_n_0 ,\shift_array[1][7]_i_9_n_0 }),
        .O(data0[7:0]),
        .S({\shift_array[1][7]_i_10_n_0 ,\shift_array[1][7]_i_11_n_0 ,\shift_array[1][7]_i_12_n_0 ,\shift_array[1][7]_i_13_n_0 ,\shift_array[1][7]_i_14_n_0 ,\shift_array[1][7]_i_15_n_0 ,\shift_array[1][7]_i_16_n_0 ,\shift_array[1][7]_i_17_n_0 }));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[8]),
        .Q(\shift_array_reg_n_0_[1][8] ),
        .R(calc_is_zero));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[9]),
        .Q(\shift_array_reg_n_0_[1][9] ),
        .R(calc_is_zero));
endmodule

(* ORIG_REF_NAME = "shiftreg" *) 
module ponos_shiftreg__parameterized1
   (calc_bucket_set_addr_i_dld,
    \gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[1][0] ,
    \DELAY_BLOCK[3].shift_array_reg[4][1]_0 ,
    \DELAY_BLOCK[3].shift_array_reg[4][1]_1 ,
    \DELAY_BLOCK[3].shift_array_reg[4][0]_0 ,
    \DELAY_BLOCK[3].shift_array_reg[4][2]_0 ,
    \DELAY_BLOCK[3].shift_array_reg[4][2]_1 ,
    \DELAY_BLOCK[3].shift_array_reg[4][0]_1 ,
    prsi_index_i,
    clk,
    douta,
    calc_is_zero_dld,
    accept_flags_o,
    calc_is_dummy_dld,
    processing_first_accept_flag,
    Q,
    \accept_flags_o_reg[2] );
  output [2:0]calc_bucket_set_addr_i_dld;
  output \gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[1][0] ;
  output \DELAY_BLOCK[3].shift_array_reg[4][1]_0 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][1]_1 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][0]_0 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][2]_0 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][2]_1 ;
  output \DELAY_BLOCK[3].shift_array_reg[4][0]_1 ;
  input [2:0]prsi_index_i;
  input clk;
  input [0:0]douta;
  input calc_is_zero_dld;
  input [2:0]accept_flags_o;
  input calc_is_dummy_dld;
  input processing_first_accept_flag;
  input [0:0]Q;
  input \accept_flags_o_reg[2] ;

  wire \<const0> ;
  wire \<const1> ;
  wire \DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ;
  wire \DELAY_BLOCK[2].shift_array_reg[3][1]_srl3_n_0 ;
  wire \DELAY_BLOCK[2].shift_array_reg[3][2]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][0]_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][0]_1 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1]_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1]_1 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][2]_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][2]_1 ;
  wire [0:0]Q;
  wire [2:0]accept_flags_o;
  wire \accept_flags_o[0]_i_2_n_0 ;
  wire \accept_flags_o[2]_i_2_n_0 ;
  wire \accept_flags_o[2]_i_3_n_0 ;
  wire \accept_flags_o[5]_i_2_n_0 ;
  wire \accept_flags_o[5]_i_3_n_0 ;
  wire \accept_flags_o_reg[2] ;
  wire [2:0]calc_bucket_set_addr_i_dld;
  wire calc_is_dummy_dld;
  wire calc_is_zero_dld;
  wire clk;
  wire [0:0]douta;
  wire \gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[1][0] ;
  wire processing_first_accept_flag;
  wire [2:0]prsi_index_i;

  (* srl_bus_name = "\\i_shiftreg_calc_bucket_set_addr/DELAY_BLOCK[2].shift_array_reg[3] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_set_addr/DELAY_BLOCK[2].shift_array_reg[3][0]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[2].shift_array_reg[3][0]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(prsi_index_i[0]),
        .Q(\DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_set_addr/DELAY_BLOCK[2].shift_array_reg[3] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_set_addr/DELAY_BLOCK[2].shift_array_reg[3][1]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[2].shift_array_reg[3][1]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(prsi_index_i[1]),
        .Q(\DELAY_BLOCK[2].shift_array_reg[3][1]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_calc_bucket_set_addr/DELAY_BLOCK[2].shift_array_reg[3] " *) 
  (* srl_name = "\\i_shiftreg_calc_bucket_set_addr/DELAY_BLOCK[2].shift_array_reg[3][2]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[2].shift_array_reg[3][2]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(prsi_index_i[2]),
        .Q(\DELAY_BLOCK[2].shift_array_reg[3][2]_srl3_n_0 ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[3].shift_array_reg[4][0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[2].shift_array_reg[3][0]_srl3_n_0 ),
        .Q(calc_bucket_set_addr_i_dld[0]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[2].shift_array_reg[3][1]_srl3_n_0 ),
        .Q(calc_bucket_set_addr_i_dld[1]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[3].shift_array_reg[4][2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[2].shift_array_reg[3][2]_srl3_n_0 ),
        .Q(calc_bucket_set_addr_i_dld[2]),
        .R(\<const0> ));
  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT6 #(
    .INIT(64'hFFFFFBFFFFFF0800)) 
    \accept_flags_o[0]_i_1 
       (.I0(\accept_flags_o_reg[2] ),
        .I1(\accept_flags_o[2]_i_2_n_0 ),
        .I2(calc_bucket_set_addr_i_dld[1]),
        .I3(Q),
        .I4(\accept_flags_o[0]_i_2_n_0 ),
        .I5(accept_flags_o[0]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][1]_1 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88888880)) 
    \accept_flags_o[0]_i_2 
       (.I0(Q),
        .I1(processing_first_accept_flag),
        .I2(calc_bucket_set_addr_i_dld[2]),
        .I3(calc_bucket_set_addr_i_dld[0]),
        .I4(calc_bucket_set_addr_i_dld[1]),
        .I5(calc_is_dummy_dld),
        .O(\accept_flags_o[0]_i_2_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \accept_flags_o[1]_i_2 
       (.I0(calc_bucket_set_addr_i_dld[0]),
        .I1(calc_bucket_set_addr_i_dld[2]),
        .I2(calc_bucket_set_addr_i_dld[1]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][0]_1 ));
  LUT6 #(
    .INIT(64'hFFFFBFFFFFFF8000)) 
    \accept_flags_o[2]_i_1 
       (.I0(\accept_flags_o_reg[2] ),
        .I1(calc_bucket_set_addr_i_dld[1]),
        .I2(\accept_flags_o[2]_i_2_n_0 ),
        .I3(Q),
        .I4(\accept_flags_o[2]_i_3_n_0 ),
        .I5(accept_flags_o[1]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][1]_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \accept_flags_o[2]_i_2 
       (.I0(calc_bucket_set_addr_i_dld[0]),
        .I1(calc_bucket_set_addr_i_dld[2]),
        .O(\accept_flags_o[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88808888)) 
    \accept_flags_o[2]_i_3 
       (.I0(Q),
        .I1(processing_first_accept_flag),
        .I2(calc_bucket_set_addr_i_dld[2]),
        .I3(calc_bucket_set_addr_i_dld[0]),
        .I4(calc_bucket_set_addr_i_dld[1]),
        .I5(calc_is_dummy_dld),
        .O(\accept_flags_o[2]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \accept_flags_o[3]_i_2 
       (.I0(calc_bucket_set_addr_i_dld[2]),
        .I1(calc_bucket_set_addr_i_dld[0]),
        .I2(calc_bucket_set_addr_i_dld[1]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][2]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \accept_flags_o[4]_i_2 
       (.I0(calc_bucket_set_addr_i_dld[2]),
        .I1(calc_bucket_set_addr_i_dld[0]),
        .I2(calc_bucket_set_addr_i_dld[1]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][2]_0 ));
  LUT5 #(
    .INIT(32'hFDFFFD00)) 
    \accept_flags_o[5]_i_1 
       (.I0(douta),
        .I1(calc_is_zero_dld),
        .I2(\accept_flags_o[5]_i_2_n_0 ),
        .I3(\accept_flags_o[5]_i_3_n_0 ),
        .I4(accept_flags_o[2]),
        .O(\gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[1][0] ));
  LUT6 #(
    .INIT(64'hAAAAAAAA88880888)) 
    \accept_flags_o[5]_i_2 
       (.I0(Q),
        .I1(processing_first_accept_flag),
        .I2(calc_bucket_set_addr_i_dld[0]),
        .I3(calc_bucket_set_addr_i_dld[2]),
        .I4(calc_bucket_set_addr_i_dld[1]),
        .I5(calc_is_dummy_dld),
        .O(\accept_flags_o[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBAAA00000000)) 
    \accept_flags_o[5]_i_3 
       (.I0(calc_is_dummy_dld),
        .I1(calc_bucket_set_addr_i_dld[1]),
        .I2(calc_bucket_set_addr_i_dld[2]),
        .I3(calc_bucket_set_addr_i_dld[0]),
        .I4(processing_first_accept_flag),
        .I5(Q),
        .O(\accept_flags_o[5]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \accept_flags_o[6]_i_3 
       (.I0(calc_bucket_set_addr_i_dld[0]),
        .I1(calc_bucket_set_addr_i_dld[2]),
        .I2(calc_bucket_set_addr_i_dld[1]),
        .O(\DELAY_BLOCK[3].shift_array_reg[4][0]_0 ));
endmodule

(* ORIG_REF_NAME = "shiftreg" *) 
module ponos_shiftreg__parameterized2
   (acc_point_o,
    clk,
    prsi_point_i);
  output [1163:0]acc_point_o;
  input clk;
  input [1163:0]prsi_point_i;

  wire \<const0> ;
  wire \<const1> ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][0]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1000]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1001]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1002]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1003]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1004]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1005]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1006]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1007]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1008]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1009]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][100]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1010]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1011]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1012]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1013]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1014]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1015]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1016]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1017]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1018]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1019]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][101]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1020]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1021]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1022]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1023]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1024]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1025]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1026]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1027]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1028]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1029]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][102]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1030]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1031]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1032]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1033]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1034]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1035]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1036]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1037]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1038]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1039]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][103]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1040]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1041]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1042]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1043]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1044]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1045]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1046]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1047]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1048]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1049]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][104]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1050]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1051]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1052]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1053]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1054]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1055]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1056]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1057]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1058]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1059]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][105]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1060]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1061]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1062]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1063]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1064]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1065]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1066]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1067]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1068]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1069]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][106]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1070]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1071]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1072]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1073]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1074]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1075]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1076]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1077]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1078]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1079]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][107]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1080]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1081]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1082]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1083]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1084]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1085]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1086]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1087]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1088]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1089]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][108]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1090]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1091]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1092]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1093]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1094]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1095]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1096]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1097]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1098]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1099]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][109]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][10]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1100]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1101]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1102]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1103]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1104]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1105]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1106]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1107]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1108]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1109]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][110]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1110]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1111]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1112]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1113]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1114]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1115]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1116]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1117]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1118]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1119]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][111]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1120]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1121]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1122]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1123]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1124]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1125]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1126]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1127]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1128]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1129]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][112]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1130]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1131]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1132]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1133]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1134]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1135]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1136]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1137]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1138]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1139]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][113]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1140]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1141]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1142]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1143]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1144]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1145]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1146]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1147]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1148]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1149]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][114]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1150]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1151]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1152]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1153]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1154]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1155]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1156]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1157]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1158]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1159]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][115]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1160]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1161]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1162]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1163]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][116]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][117]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][118]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][119]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][11]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][120]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][121]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][122]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][123]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][124]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][125]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][126]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][127]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][128]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][129]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][12]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][130]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][131]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][132]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][133]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][134]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][135]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][136]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][137]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][138]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][139]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][13]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][140]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][141]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][142]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][143]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][144]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][145]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][146]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][147]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][148]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][149]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][14]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][150]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][151]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][152]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][153]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][154]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][155]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][156]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][157]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][158]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][159]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][15]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][160]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][161]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][162]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][163]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][164]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][165]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][166]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][167]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][168]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][169]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][16]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][170]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][171]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][172]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][173]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][174]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][175]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][176]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][177]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][178]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][179]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][17]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][180]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][181]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][182]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][183]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][184]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][185]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][186]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][187]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][188]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][189]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][18]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][190]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][191]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][192]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][193]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][194]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][195]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][196]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][197]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][198]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][199]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][19]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][1]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][200]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][201]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][202]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][203]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][204]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][205]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][206]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][207]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][208]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][209]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][20]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][210]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][211]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][212]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][213]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][214]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][215]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][216]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][217]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][218]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][219]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][21]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][220]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][221]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][222]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][223]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][224]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][225]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][226]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][227]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][228]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][229]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][22]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][230]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][231]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][232]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][233]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][234]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][235]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][236]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][237]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][238]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][239]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][23]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][240]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][241]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][242]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][243]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][244]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][245]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][246]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][247]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][248]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][249]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][24]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][250]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][251]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][252]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][253]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][254]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][255]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][256]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][257]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][258]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][259]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][25]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][260]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][261]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][262]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][263]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][264]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][265]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][266]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][267]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][268]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][269]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][26]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][270]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][271]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][272]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][273]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][274]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][275]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][276]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][277]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][278]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][279]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][27]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][280]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][281]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][282]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][283]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][284]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][285]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][286]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][287]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][288]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][289]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][28]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][290]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][291]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][292]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][293]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][294]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][295]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][296]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][297]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][298]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][299]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][29]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][2]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][300]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][301]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][302]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][303]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][304]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][305]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][306]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][307]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][308]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][309]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][30]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][310]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][311]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][312]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][313]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][314]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][315]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][316]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][317]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][318]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][319]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][31]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][320]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][321]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][322]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][323]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][324]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][325]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][326]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][327]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][328]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][329]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][32]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][330]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][331]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][332]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][333]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][334]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][335]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][336]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][337]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][338]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][339]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][33]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][340]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][341]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][342]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][343]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][344]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][345]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][346]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][347]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][348]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][349]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][34]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][350]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][351]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][352]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][353]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][354]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][355]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][356]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][357]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][358]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][359]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][35]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][360]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][361]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][362]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][363]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][364]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][365]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][366]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][367]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][368]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][369]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][36]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][370]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][371]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][372]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][373]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][374]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][375]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][376]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][377]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][378]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][379]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][37]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][380]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][381]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][382]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][383]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][384]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][385]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][386]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][387]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][388]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][389]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][38]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][390]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][391]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][392]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][393]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][394]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][395]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][396]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][397]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][398]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][399]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][39]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][3]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][400]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][401]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][402]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][403]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][404]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][405]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][406]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][407]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][408]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][409]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][40]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][410]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][411]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][412]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][413]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][414]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][415]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][416]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][417]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][418]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][419]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][41]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][420]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][421]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][422]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][423]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][424]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][425]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][426]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][427]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][428]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][429]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][42]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][430]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][431]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][432]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][433]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][434]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][435]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][436]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][437]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][438]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][439]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][43]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][440]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][441]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][442]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][443]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][444]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][445]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][446]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][447]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][448]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][449]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][44]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][450]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][451]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][452]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][453]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][454]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][455]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][456]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][457]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][458]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][459]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][45]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][460]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][461]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][462]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][463]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][464]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][465]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][466]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][467]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][468]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][469]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][46]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][470]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][471]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][472]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][473]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][474]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][475]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][476]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][477]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][478]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][479]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][47]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][480]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][481]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][482]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][483]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][484]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][485]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][486]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][487]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][488]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][489]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][48]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][490]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][491]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][492]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][493]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][494]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][495]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][496]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][497]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][498]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][499]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][49]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][4]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][500]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][501]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][502]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][503]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][504]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][505]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][506]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][507]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][508]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][509]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][50]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][510]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][511]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][512]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][513]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][514]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][515]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][516]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][517]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][518]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][519]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][51]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][520]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][521]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][522]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][523]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][524]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][525]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][526]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][527]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][528]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][529]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][52]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][530]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][531]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][532]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][533]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][534]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][535]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][536]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][537]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][538]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][539]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][53]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][540]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][541]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][542]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][543]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][544]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][545]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][546]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][547]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][548]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][549]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][54]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][550]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][551]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][552]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][553]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][554]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][555]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][556]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][557]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][558]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][559]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][55]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][560]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][561]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][562]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][563]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][564]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][565]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][566]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][567]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][568]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][569]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][56]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][570]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][571]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][572]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][573]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][574]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][575]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][576]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][577]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][578]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][579]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][57]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][580]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][581]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][582]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][583]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][584]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][585]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][586]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][587]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][588]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][589]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][58]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][590]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][591]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][592]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][593]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][594]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][595]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][596]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][597]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][598]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][599]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][59]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][5]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][600]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][601]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][602]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][603]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][604]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][605]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][606]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][607]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][608]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][609]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][60]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][610]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][611]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][612]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][613]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][614]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][615]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][616]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][617]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][618]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][619]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][61]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][620]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][621]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][622]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][623]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][624]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][625]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][626]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][627]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][628]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][629]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][62]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][630]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][631]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][632]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][633]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][634]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][635]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][636]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][637]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][638]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][639]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][63]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][640]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][641]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][642]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][643]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][644]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][645]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][646]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][647]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][648]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][649]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][64]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][650]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][651]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][652]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][653]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][654]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][655]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][656]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][657]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][658]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][659]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][65]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][660]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][661]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][662]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][663]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][664]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][665]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][666]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][667]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][668]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][669]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][66]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][670]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][671]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][672]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][673]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][674]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][675]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][676]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][677]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][678]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][679]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][67]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][680]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][681]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][682]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][683]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][684]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][685]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][686]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][687]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][688]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][689]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][68]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][690]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][691]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][692]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][693]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][694]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][695]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][696]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][697]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][698]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][699]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][69]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][6]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][700]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][701]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][702]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][703]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][704]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][705]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][706]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][707]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][708]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][709]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][70]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][710]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][711]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][712]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][713]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][714]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][715]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][716]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][717]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][718]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][719]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][71]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][720]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][721]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][722]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][723]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][724]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][725]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][726]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][727]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][728]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][729]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][72]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][730]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][731]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][732]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][733]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][734]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][735]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][736]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][737]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][738]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][739]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][73]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][740]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][741]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][742]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][743]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][744]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][745]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][746]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][747]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][748]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][749]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][74]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][750]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][751]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][752]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][753]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][754]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][755]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][756]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][757]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][758]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][759]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][75]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][760]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][761]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][762]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][763]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][764]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][765]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][766]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][767]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][768]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][769]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][76]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][770]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][771]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][772]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][773]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][774]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][775]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][776]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][777]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][778]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][779]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][77]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][780]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][781]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][782]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][783]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][784]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][785]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][786]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][787]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][788]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][789]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][78]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][790]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][791]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][792]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][793]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][794]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][795]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][796]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][797]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][798]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][799]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][79]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][7]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][800]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][801]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][802]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][803]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][804]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][805]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][806]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][807]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][808]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][809]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][80]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][810]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][811]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][812]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][813]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][814]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][815]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][816]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][817]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][818]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][819]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][81]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][820]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][821]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][822]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][823]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][824]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][825]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][826]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][827]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][828]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][829]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][82]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][830]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][831]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][832]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][833]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][834]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][835]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][836]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][837]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][838]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][839]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][83]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][840]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][841]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][842]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][843]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][844]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][845]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][846]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][847]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][848]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][849]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][84]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][850]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][851]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][852]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][853]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][854]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][855]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][856]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][857]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][858]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][859]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][85]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][860]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][861]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][862]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][863]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][864]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][865]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][866]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][867]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][868]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][869]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][86]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][870]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][871]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][872]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][873]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][874]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][875]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][876]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][877]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][878]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][879]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][87]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][880]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][881]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][882]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][883]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][884]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][885]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][886]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][887]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][888]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][889]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][88]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][890]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][891]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][892]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][893]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][894]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][895]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][896]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][897]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][898]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][899]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][89]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][8]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][900]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][901]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][902]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][903]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][904]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][905]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][906]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][907]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][908]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][909]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][90]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][910]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][911]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][912]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][913]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][914]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][915]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][916]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][917]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][918]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][919]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][91]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][920]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][921]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][922]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][923]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][924]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][925]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][926]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][927]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][928]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][929]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][92]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][930]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][931]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][932]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][933]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][934]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][935]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][936]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][937]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][938]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][939]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][93]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][940]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][941]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][942]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][943]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][944]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][945]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][946]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][947]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][948]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][949]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][94]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][950]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][951]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][952]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][953]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][954]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][955]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][956]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][957]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][958]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][959]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][95]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][960]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][961]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][962]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][963]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][964]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][965]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][966]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][967]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][968]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][969]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][96]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][970]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][971]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][972]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][973]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][974]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][975]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][976]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][977]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][978]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][979]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][97]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][980]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][981]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][982]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][983]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][984]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][985]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][986]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][987]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][988]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][989]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][98]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][990]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][991]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][992]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][993]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][994]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][995]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][996]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][997]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][998]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][999]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][99]_srl3_n_0 ;
  wire \DELAY_BLOCK[3].shift_array_reg[4][9]_srl3_n_0 ;
  wire [1163:0]acc_point_o;
  wire clk;
  wire [1163:0]prsi_point_i;
  wire \shift_array_reg_n_0_[1][0] ;
  wire \shift_array_reg_n_0_[1][1000] ;
  wire \shift_array_reg_n_0_[1][1001] ;
  wire \shift_array_reg_n_0_[1][1002] ;
  wire \shift_array_reg_n_0_[1][1003] ;
  wire \shift_array_reg_n_0_[1][1004] ;
  wire \shift_array_reg_n_0_[1][1005] ;
  wire \shift_array_reg_n_0_[1][1006] ;
  wire \shift_array_reg_n_0_[1][1007] ;
  wire \shift_array_reg_n_0_[1][1008] ;
  wire \shift_array_reg_n_0_[1][1009] ;
  wire \shift_array_reg_n_0_[1][100] ;
  wire \shift_array_reg_n_0_[1][1010] ;
  wire \shift_array_reg_n_0_[1][1011] ;
  wire \shift_array_reg_n_0_[1][1012] ;
  wire \shift_array_reg_n_0_[1][1013] ;
  wire \shift_array_reg_n_0_[1][1014] ;
  wire \shift_array_reg_n_0_[1][1015] ;
  wire \shift_array_reg_n_0_[1][1016] ;
  wire \shift_array_reg_n_0_[1][1017] ;
  wire \shift_array_reg_n_0_[1][1018] ;
  wire \shift_array_reg_n_0_[1][1019] ;
  wire \shift_array_reg_n_0_[1][101] ;
  wire \shift_array_reg_n_0_[1][1020] ;
  wire \shift_array_reg_n_0_[1][1021] ;
  wire \shift_array_reg_n_0_[1][1022] ;
  wire \shift_array_reg_n_0_[1][1023] ;
  wire \shift_array_reg_n_0_[1][1024] ;
  wire \shift_array_reg_n_0_[1][1025] ;
  wire \shift_array_reg_n_0_[1][1026] ;
  wire \shift_array_reg_n_0_[1][1027] ;
  wire \shift_array_reg_n_0_[1][1028] ;
  wire \shift_array_reg_n_0_[1][1029] ;
  wire \shift_array_reg_n_0_[1][102] ;
  wire \shift_array_reg_n_0_[1][1030] ;
  wire \shift_array_reg_n_0_[1][1031] ;
  wire \shift_array_reg_n_0_[1][1032] ;
  wire \shift_array_reg_n_0_[1][1033] ;
  wire \shift_array_reg_n_0_[1][1034] ;
  wire \shift_array_reg_n_0_[1][1035] ;
  wire \shift_array_reg_n_0_[1][1036] ;
  wire \shift_array_reg_n_0_[1][1037] ;
  wire \shift_array_reg_n_0_[1][1038] ;
  wire \shift_array_reg_n_0_[1][1039] ;
  wire \shift_array_reg_n_0_[1][103] ;
  wire \shift_array_reg_n_0_[1][1040] ;
  wire \shift_array_reg_n_0_[1][1041] ;
  wire \shift_array_reg_n_0_[1][1042] ;
  wire \shift_array_reg_n_0_[1][1043] ;
  wire \shift_array_reg_n_0_[1][1044] ;
  wire \shift_array_reg_n_0_[1][1045] ;
  wire \shift_array_reg_n_0_[1][1046] ;
  wire \shift_array_reg_n_0_[1][1047] ;
  wire \shift_array_reg_n_0_[1][1048] ;
  wire \shift_array_reg_n_0_[1][1049] ;
  wire \shift_array_reg_n_0_[1][104] ;
  wire \shift_array_reg_n_0_[1][1050] ;
  wire \shift_array_reg_n_0_[1][1051] ;
  wire \shift_array_reg_n_0_[1][1052] ;
  wire \shift_array_reg_n_0_[1][1053] ;
  wire \shift_array_reg_n_0_[1][1054] ;
  wire \shift_array_reg_n_0_[1][1055] ;
  wire \shift_array_reg_n_0_[1][1056] ;
  wire \shift_array_reg_n_0_[1][1057] ;
  wire \shift_array_reg_n_0_[1][1058] ;
  wire \shift_array_reg_n_0_[1][1059] ;
  wire \shift_array_reg_n_0_[1][105] ;
  wire \shift_array_reg_n_0_[1][1060] ;
  wire \shift_array_reg_n_0_[1][1061] ;
  wire \shift_array_reg_n_0_[1][1062] ;
  wire \shift_array_reg_n_0_[1][1063] ;
  wire \shift_array_reg_n_0_[1][1064] ;
  wire \shift_array_reg_n_0_[1][1065] ;
  wire \shift_array_reg_n_0_[1][1066] ;
  wire \shift_array_reg_n_0_[1][1067] ;
  wire \shift_array_reg_n_0_[1][1068] ;
  wire \shift_array_reg_n_0_[1][1069] ;
  wire \shift_array_reg_n_0_[1][106] ;
  wire \shift_array_reg_n_0_[1][1070] ;
  wire \shift_array_reg_n_0_[1][1071] ;
  wire \shift_array_reg_n_0_[1][1072] ;
  wire \shift_array_reg_n_0_[1][1073] ;
  wire \shift_array_reg_n_0_[1][1074] ;
  wire \shift_array_reg_n_0_[1][1075] ;
  wire \shift_array_reg_n_0_[1][1076] ;
  wire \shift_array_reg_n_0_[1][1077] ;
  wire \shift_array_reg_n_0_[1][1078] ;
  wire \shift_array_reg_n_0_[1][1079] ;
  wire \shift_array_reg_n_0_[1][107] ;
  wire \shift_array_reg_n_0_[1][1080] ;
  wire \shift_array_reg_n_0_[1][1081] ;
  wire \shift_array_reg_n_0_[1][1082] ;
  wire \shift_array_reg_n_0_[1][1083] ;
  wire \shift_array_reg_n_0_[1][1084] ;
  wire \shift_array_reg_n_0_[1][1085] ;
  wire \shift_array_reg_n_0_[1][1086] ;
  wire \shift_array_reg_n_0_[1][1087] ;
  wire \shift_array_reg_n_0_[1][1088] ;
  wire \shift_array_reg_n_0_[1][1089] ;
  wire \shift_array_reg_n_0_[1][108] ;
  wire \shift_array_reg_n_0_[1][1090] ;
  wire \shift_array_reg_n_0_[1][1091] ;
  wire \shift_array_reg_n_0_[1][1092] ;
  wire \shift_array_reg_n_0_[1][1093] ;
  wire \shift_array_reg_n_0_[1][1094] ;
  wire \shift_array_reg_n_0_[1][1095] ;
  wire \shift_array_reg_n_0_[1][1096] ;
  wire \shift_array_reg_n_0_[1][1097] ;
  wire \shift_array_reg_n_0_[1][1098] ;
  wire \shift_array_reg_n_0_[1][1099] ;
  wire \shift_array_reg_n_0_[1][109] ;
  wire \shift_array_reg_n_0_[1][10] ;
  wire \shift_array_reg_n_0_[1][1100] ;
  wire \shift_array_reg_n_0_[1][1101] ;
  wire \shift_array_reg_n_0_[1][1102] ;
  wire \shift_array_reg_n_0_[1][1103] ;
  wire \shift_array_reg_n_0_[1][1104] ;
  wire \shift_array_reg_n_0_[1][1105] ;
  wire \shift_array_reg_n_0_[1][1106] ;
  wire \shift_array_reg_n_0_[1][1107] ;
  wire \shift_array_reg_n_0_[1][1108] ;
  wire \shift_array_reg_n_0_[1][1109] ;
  wire \shift_array_reg_n_0_[1][110] ;
  wire \shift_array_reg_n_0_[1][1110] ;
  wire \shift_array_reg_n_0_[1][1111] ;
  wire \shift_array_reg_n_0_[1][1112] ;
  wire \shift_array_reg_n_0_[1][1113] ;
  wire \shift_array_reg_n_0_[1][1114] ;
  wire \shift_array_reg_n_0_[1][1115] ;
  wire \shift_array_reg_n_0_[1][1116] ;
  wire \shift_array_reg_n_0_[1][1117] ;
  wire \shift_array_reg_n_0_[1][1118] ;
  wire \shift_array_reg_n_0_[1][1119] ;
  wire \shift_array_reg_n_0_[1][111] ;
  wire \shift_array_reg_n_0_[1][1120] ;
  wire \shift_array_reg_n_0_[1][1121] ;
  wire \shift_array_reg_n_0_[1][1122] ;
  wire \shift_array_reg_n_0_[1][1123] ;
  wire \shift_array_reg_n_0_[1][1124] ;
  wire \shift_array_reg_n_0_[1][1125] ;
  wire \shift_array_reg_n_0_[1][1126] ;
  wire \shift_array_reg_n_0_[1][1127] ;
  wire \shift_array_reg_n_0_[1][1128] ;
  wire \shift_array_reg_n_0_[1][1129] ;
  wire \shift_array_reg_n_0_[1][112] ;
  wire \shift_array_reg_n_0_[1][1130] ;
  wire \shift_array_reg_n_0_[1][1131] ;
  wire \shift_array_reg_n_0_[1][1132] ;
  wire \shift_array_reg_n_0_[1][1133] ;
  wire \shift_array_reg_n_0_[1][1134] ;
  wire \shift_array_reg_n_0_[1][1135] ;
  wire \shift_array_reg_n_0_[1][1136] ;
  wire \shift_array_reg_n_0_[1][1137] ;
  wire \shift_array_reg_n_0_[1][1138] ;
  wire \shift_array_reg_n_0_[1][1139] ;
  wire \shift_array_reg_n_0_[1][113] ;
  wire \shift_array_reg_n_0_[1][1140] ;
  wire \shift_array_reg_n_0_[1][1141] ;
  wire \shift_array_reg_n_0_[1][1142] ;
  wire \shift_array_reg_n_0_[1][1143] ;
  wire \shift_array_reg_n_0_[1][1144] ;
  wire \shift_array_reg_n_0_[1][1145] ;
  wire \shift_array_reg_n_0_[1][1146] ;
  wire \shift_array_reg_n_0_[1][1147] ;
  wire \shift_array_reg_n_0_[1][1148] ;
  wire \shift_array_reg_n_0_[1][1149] ;
  wire \shift_array_reg_n_0_[1][114] ;
  wire \shift_array_reg_n_0_[1][1150] ;
  wire \shift_array_reg_n_0_[1][1151] ;
  wire \shift_array_reg_n_0_[1][1152] ;
  wire \shift_array_reg_n_0_[1][1153] ;
  wire \shift_array_reg_n_0_[1][1154] ;
  wire \shift_array_reg_n_0_[1][1155] ;
  wire \shift_array_reg_n_0_[1][1156] ;
  wire \shift_array_reg_n_0_[1][1157] ;
  wire \shift_array_reg_n_0_[1][1158] ;
  wire \shift_array_reg_n_0_[1][1159] ;
  wire \shift_array_reg_n_0_[1][115] ;
  wire \shift_array_reg_n_0_[1][1160] ;
  wire \shift_array_reg_n_0_[1][1161] ;
  wire \shift_array_reg_n_0_[1][1162] ;
  wire \shift_array_reg_n_0_[1][1163] ;
  wire \shift_array_reg_n_0_[1][116] ;
  wire \shift_array_reg_n_0_[1][117] ;
  wire \shift_array_reg_n_0_[1][118] ;
  wire \shift_array_reg_n_0_[1][119] ;
  wire \shift_array_reg_n_0_[1][11] ;
  wire \shift_array_reg_n_0_[1][120] ;
  wire \shift_array_reg_n_0_[1][121] ;
  wire \shift_array_reg_n_0_[1][122] ;
  wire \shift_array_reg_n_0_[1][123] ;
  wire \shift_array_reg_n_0_[1][124] ;
  wire \shift_array_reg_n_0_[1][125] ;
  wire \shift_array_reg_n_0_[1][126] ;
  wire \shift_array_reg_n_0_[1][127] ;
  wire \shift_array_reg_n_0_[1][128] ;
  wire \shift_array_reg_n_0_[1][129] ;
  wire \shift_array_reg_n_0_[1][12] ;
  wire \shift_array_reg_n_0_[1][130] ;
  wire \shift_array_reg_n_0_[1][131] ;
  wire \shift_array_reg_n_0_[1][132] ;
  wire \shift_array_reg_n_0_[1][133] ;
  wire \shift_array_reg_n_0_[1][134] ;
  wire \shift_array_reg_n_0_[1][135] ;
  wire \shift_array_reg_n_0_[1][136] ;
  wire \shift_array_reg_n_0_[1][137] ;
  wire \shift_array_reg_n_0_[1][138] ;
  wire \shift_array_reg_n_0_[1][139] ;
  wire \shift_array_reg_n_0_[1][13] ;
  wire \shift_array_reg_n_0_[1][140] ;
  wire \shift_array_reg_n_0_[1][141] ;
  wire \shift_array_reg_n_0_[1][142] ;
  wire \shift_array_reg_n_0_[1][143] ;
  wire \shift_array_reg_n_0_[1][144] ;
  wire \shift_array_reg_n_0_[1][145] ;
  wire \shift_array_reg_n_0_[1][146] ;
  wire \shift_array_reg_n_0_[1][147] ;
  wire \shift_array_reg_n_0_[1][148] ;
  wire \shift_array_reg_n_0_[1][149] ;
  wire \shift_array_reg_n_0_[1][14] ;
  wire \shift_array_reg_n_0_[1][150] ;
  wire \shift_array_reg_n_0_[1][151] ;
  wire \shift_array_reg_n_0_[1][152] ;
  wire \shift_array_reg_n_0_[1][153] ;
  wire \shift_array_reg_n_0_[1][154] ;
  wire \shift_array_reg_n_0_[1][155] ;
  wire \shift_array_reg_n_0_[1][156] ;
  wire \shift_array_reg_n_0_[1][157] ;
  wire \shift_array_reg_n_0_[1][158] ;
  wire \shift_array_reg_n_0_[1][159] ;
  wire \shift_array_reg_n_0_[1][15] ;
  wire \shift_array_reg_n_0_[1][160] ;
  wire \shift_array_reg_n_0_[1][161] ;
  wire \shift_array_reg_n_0_[1][162] ;
  wire \shift_array_reg_n_0_[1][163] ;
  wire \shift_array_reg_n_0_[1][164] ;
  wire \shift_array_reg_n_0_[1][165] ;
  wire \shift_array_reg_n_0_[1][166] ;
  wire \shift_array_reg_n_0_[1][167] ;
  wire \shift_array_reg_n_0_[1][168] ;
  wire \shift_array_reg_n_0_[1][169] ;
  wire \shift_array_reg_n_0_[1][16] ;
  wire \shift_array_reg_n_0_[1][170] ;
  wire \shift_array_reg_n_0_[1][171] ;
  wire \shift_array_reg_n_0_[1][172] ;
  wire \shift_array_reg_n_0_[1][173] ;
  wire \shift_array_reg_n_0_[1][174] ;
  wire \shift_array_reg_n_0_[1][175] ;
  wire \shift_array_reg_n_0_[1][176] ;
  wire \shift_array_reg_n_0_[1][177] ;
  wire \shift_array_reg_n_0_[1][178] ;
  wire \shift_array_reg_n_0_[1][179] ;
  wire \shift_array_reg_n_0_[1][17] ;
  wire \shift_array_reg_n_0_[1][180] ;
  wire \shift_array_reg_n_0_[1][181] ;
  wire \shift_array_reg_n_0_[1][182] ;
  wire \shift_array_reg_n_0_[1][183] ;
  wire \shift_array_reg_n_0_[1][184] ;
  wire \shift_array_reg_n_0_[1][185] ;
  wire \shift_array_reg_n_0_[1][186] ;
  wire \shift_array_reg_n_0_[1][187] ;
  wire \shift_array_reg_n_0_[1][188] ;
  wire \shift_array_reg_n_0_[1][189] ;
  wire \shift_array_reg_n_0_[1][18] ;
  wire \shift_array_reg_n_0_[1][190] ;
  wire \shift_array_reg_n_0_[1][191] ;
  wire \shift_array_reg_n_0_[1][192] ;
  wire \shift_array_reg_n_0_[1][193] ;
  wire \shift_array_reg_n_0_[1][194] ;
  wire \shift_array_reg_n_0_[1][195] ;
  wire \shift_array_reg_n_0_[1][196] ;
  wire \shift_array_reg_n_0_[1][197] ;
  wire \shift_array_reg_n_0_[1][198] ;
  wire \shift_array_reg_n_0_[1][199] ;
  wire \shift_array_reg_n_0_[1][19] ;
  wire \shift_array_reg_n_0_[1][1] ;
  wire \shift_array_reg_n_0_[1][200] ;
  wire \shift_array_reg_n_0_[1][201] ;
  wire \shift_array_reg_n_0_[1][202] ;
  wire \shift_array_reg_n_0_[1][203] ;
  wire \shift_array_reg_n_0_[1][204] ;
  wire \shift_array_reg_n_0_[1][205] ;
  wire \shift_array_reg_n_0_[1][206] ;
  wire \shift_array_reg_n_0_[1][207] ;
  wire \shift_array_reg_n_0_[1][208] ;
  wire \shift_array_reg_n_0_[1][209] ;
  wire \shift_array_reg_n_0_[1][20] ;
  wire \shift_array_reg_n_0_[1][210] ;
  wire \shift_array_reg_n_0_[1][211] ;
  wire \shift_array_reg_n_0_[1][212] ;
  wire \shift_array_reg_n_0_[1][213] ;
  wire \shift_array_reg_n_0_[1][214] ;
  wire \shift_array_reg_n_0_[1][215] ;
  wire \shift_array_reg_n_0_[1][216] ;
  wire \shift_array_reg_n_0_[1][217] ;
  wire \shift_array_reg_n_0_[1][218] ;
  wire \shift_array_reg_n_0_[1][219] ;
  wire \shift_array_reg_n_0_[1][21] ;
  wire \shift_array_reg_n_0_[1][220] ;
  wire \shift_array_reg_n_0_[1][221] ;
  wire \shift_array_reg_n_0_[1][222] ;
  wire \shift_array_reg_n_0_[1][223] ;
  wire \shift_array_reg_n_0_[1][224] ;
  wire \shift_array_reg_n_0_[1][225] ;
  wire \shift_array_reg_n_0_[1][226] ;
  wire \shift_array_reg_n_0_[1][227] ;
  wire \shift_array_reg_n_0_[1][228] ;
  wire \shift_array_reg_n_0_[1][229] ;
  wire \shift_array_reg_n_0_[1][22] ;
  wire \shift_array_reg_n_0_[1][230] ;
  wire \shift_array_reg_n_0_[1][231] ;
  wire \shift_array_reg_n_0_[1][232] ;
  wire \shift_array_reg_n_0_[1][233] ;
  wire \shift_array_reg_n_0_[1][234] ;
  wire \shift_array_reg_n_0_[1][235] ;
  wire \shift_array_reg_n_0_[1][236] ;
  wire \shift_array_reg_n_0_[1][237] ;
  wire \shift_array_reg_n_0_[1][238] ;
  wire \shift_array_reg_n_0_[1][239] ;
  wire \shift_array_reg_n_0_[1][23] ;
  wire \shift_array_reg_n_0_[1][240] ;
  wire \shift_array_reg_n_0_[1][241] ;
  wire \shift_array_reg_n_0_[1][242] ;
  wire \shift_array_reg_n_0_[1][243] ;
  wire \shift_array_reg_n_0_[1][244] ;
  wire \shift_array_reg_n_0_[1][245] ;
  wire \shift_array_reg_n_0_[1][246] ;
  wire \shift_array_reg_n_0_[1][247] ;
  wire \shift_array_reg_n_0_[1][248] ;
  wire \shift_array_reg_n_0_[1][249] ;
  wire \shift_array_reg_n_0_[1][24] ;
  wire \shift_array_reg_n_0_[1][250] ;
  wire \shift_array_reg_n_0_[1][251] ;
  wire \shift_array_reg_n_0_[1][252] ;
  wire \shift_array_reg_n_0_[1][253] ;
  wire \shift_array_reg_n_0_[1][254] ;
  wire \shift_array_reg_n_0_[1][255] ;
  wire \shift_array_reg_n_0_[1][256] ;
  wire \shift_array_reg_n_0_[1][257] ;
  wire \shift_array_reg_n_0_[1][258] ;
  wire \shift_array_reg_n_0_[1][259] ;
  wire \shift_array_reg_n_0_[1][25] ;
  wire \shift_array_reg_n_0_[1][260] ;
  wire \shift_array_reg_n_0_[1][261] ;
  wire \shift_array_reg_n_0_[1][262] ;
  wire \shift_array_reg_n_0_[1][263] ;
  wire \shift_array_reg_n_0_[1][264] ;
  wire \shift_array_reg_n_0_[1][265] ;
  wire \shift_array_reg_n_0_[1][266] ;
  wire \shift_array_reg_n_0_[1][267] ;
  wire \shift_array_reg_n_0_[1][268] ;
  wire \shift_array_reg_n_0_[1][269] ;
  wire \shift_array_reg_n_0_[1][26] ;
  wire \shift_array_reg_n_0_[1][270] ;
  wire \shift_array_reg_n_0_[1][271] ;
  wire \shift_array_reg_n_0_[1][272] ;
  wire \shift_array_reg_n_0_[1][273] ;
  wire \shift_array_reg_n_0_[1][274] ;
  wire \shift_array_reg_n_0_[1][275] ;
  wire \shift_array_reg_n_0_[1][276] ;
  wire \shift_array_reg_n_0_[1][277] ;
  wire \shift_array_reg_n_0_[1][278] ;
  wire \shift_array_reg_n_0_[1][279] ;
  wire \shift_array_reg_n_0_[1][27] ;
  wire \shift_array_reg_n_0_[1][280] ;
  wire \shift_array_reg_n_0_[1][281] ;
  wire \shift_array_reg_n_0_[1][282] ;
  wire \shift_array_reg_n_0_[1][283] ;
  wire \shift_array_reg_n_0_[1][284] ;
  wire \shift_array_reg_n_0_[1][285] ;
  wire \shift_array_reg_n_0_[1][286] ;
  wire \shift_array_reg_n_0_[1][287] ;
  wire \shift_array_reg_n_0_[1][288] ;
  wire \shift_array_reg_n_0_[1][289] ;
  wire \shift_array_reg_n_0_[1][28] ;
  wire \shift_array_reg_n_0_[1][290] ;
  wire \shift_array_reg_n_0_[1][291] ;
  wire \shift_array_reg_n_0_[1][292] ;
  wire \shift_array_reg_n_0_[1][293] ;
  wire \shift_array_reg_n_0_[1][294] ;
  wire \shift_array_reg_n_0_[1][295] ;
  wire \shift_array_reg_n_0_[1][296] ;
  wire \shift_array_reg_n_0_[1][297] ;
  wire \shift_array_reg_n_0_[1][298] ;
  wire \shift_array_reg_n_0_[1][299] ;
  wire \shift_array_reg_n_0_[1][29] ;
  wire \shift_array_reg_n_0_[1][2] ;
  wire \shift_array_reg_n_0_[1][300] ;
  wire \shift_array_reg_n_0_[1][301] ;
  wire \shift_array_reg_n_0_[1][302] ;
  wire \shift_array_reg_n_0_[1][303] ;
  wire \shift_array_reg_n_0_[1][304] ;
  wire \shift_array_reg_n_0_[1][305] ;
  wire \shift_array_reg_n_0_[1][306] ;
  wire \shift_array_reg_n_0_[1][307] ;
  wire \shift_array_reg_n_0_[1][308] ;
  wire \shift_array_reg_n_0_[1][309] ;
  wire \shift_array_reg_n_0_[1][30] ;
  wire \shift_array_reg_n_0_[1][310] ;
  wire \shift_array_reg_n_0_[1][311] ;
  wire \shift_array_reg_n_0_[1][312] ;
  wire \shift_array_reg_n_0_[1][313] ;
  wire \shift_array_reg_n_0_[1][314] ;
  wire \shift_array_reg_n_0_[1][315] ;
  wire \shift_array_reg_n_0_[1][316] ;
  wire \shift_array_reg_n_0_[1][317] ;
  wire \shift_array_reg_n_0_[1][318] ;
  wire \shift_array_reg_n_0_[1][319] ;
  wire \shift_array_reg_n_0_[1][31] ;
  wire \shift_array_reg_n_0_[1][320] ;
  wire \shift_array_reg_n_0_[1][321] ;
  wire \shift_array_reg_n_0_[1][322] ;
  wire \shift_array_reg_n_0_[1][323] ;
  wire \shift_array_reg_n_0_[1][324] ;
  wire \shift_array_reg_n_0_[1][325] ;
  wire \shift_array_reg_n_0_[1][326] ;
  wire \shift_array_reg_n_0_[1][327] ;
  wire \shift_array_reg_n_0_[1][328] ;
  wire \shift_array_reg_n_0_[1][329] ;
  wire \shift_array_reg_n_0_[1][32] ;
  wire \shift_array_reg_n_0_[1][330] ;
  wire \shift_array_reg_n_0_[1][331] ;
  wire \shift_array_reg_n_0_[1][332] ;
  wire \shift_array_reg_n_0_[1][333] ;
  wire \shift_array_reg_n_0_[1][334] ;
  wire \shift_array_reg_n_0_[1][335] ;
  wire \shift_array_reg_n_0_[1][336] ;
  wire \shift_array_reg_n_0_[1][337] ;
  wire \shift_array_reg_n_0_[1][338] ;
  wire \shift_array_reg_n_0_[1][339] ;
  wire \shift_array_reg_n_0_[1][33] ;
  wire \shift_array_reg_n_0_[1][340] ;
  wire \shift_array_reg_n_0_[1][341] ;
  wire \shift_array_reg_n_0_[1][342] ;
  wire \shift_array_reg_n_0_[1][343] ;
  wire \shift_array_reg_n_0_[1][344] ;
  wire \shift_array_reg_n_0_[1][345] ;
  wire \shift_array_reg_n_0_[1][346] ;
  wire \shift_array_reg_n_0_[1][347] ;
  wire \shift_array_reg_n_0_[1][348] ;
  wire \shift_array_reg_n_0_[1][349] ;
  wire \shift_array_reg_n_0_[1][34] ;
  wire \shift_array_reg_n_0_[1][350] ;
  wire \shift_array_reg_n_0_[1][351] ;
  wire \shift_array_reg_n_0_[1][352] ;
  wire \shift_array_reg_n_0_[1][353] ;
  wire \shift_array_reg_n_0_[1][354] ;
  wire \shift_array_reg_n_0_[1][355] ;
  wire \shift_array_reg_n_0_[1][356] ;
  wire \shift_array_reg_n_0_[1][357] ;
  wire \shift_array_reg_n_0_[1][358] ;
  wire \shift_array_reg_n_0_[1][359] ;
  wire \shift_array_reg_n_0_[1][35] ;
  wire \shift_array_reg_n_0_[1][360] ;
  wire \shift_array_reg_n_0_[1][361] ;
  wire \shift_array_reg_n_0_[1][362] ;
  wire \shift_array_reg_n_0_[1][363] ;
  wire \shift_array_reg_n_0_[1][364] ;
  wire \shift_array_reg_n_0_[1][365] ;
  wire \shift_array_reg_n_0_[1][366] ;
  wire \shift_array_reg_n_0_[1][367] ;
  wire \shift_array_reg_n_0_[1][368] ;
  wire \shift_array_reg_n_0_[1][369] ;
  wire \shift_array_reg_n_0_[1][36] ;
  wire \shift_array_reg_n_0_[1][370] ;
  wire \shift_array_reg_n_0_[1][371] ;
  wire \shift_array_reg_n_0_[1][372] ;
  wire \shift_array_reg_n_0_[1][373] ;
  wire \shift_array_reg_n_0_[1][374] ;
  wire \shift_array_reg_n_0_[1][375] ;
  wire \shift_array_reg_n_0_[1][376] ;
  wire \shift_array_reg_n_0_[1][377] ;
  wire \shift_array_reg_n_0_[1][378] ;
  wire \shift_array_reg_n_0_[1][379] ;
  wire \shift_array_reg_n_0_[1][37] ;
  wire \shift_array_reg_n_0_[1][380] ;
  wire \shift_array_reg_n_0_[1][381] ;
  wire \shift_array_reg_n_0_[1][382] ;
  wire \shift_array_reg_n_0_[1][383] ;
  wire \shift_array_reg_n_0_[1][384] ;
  wire \shift_array_reg_n_0_[1][385] ;
  wire \shift_array_reg_n_0_[1][386] ;
  wire \shift_array_reg_n_0_[1][387] ;
  wire \shift_array_reg_n_0_[1][388] ;
  wire \shift_array_reg_n_0_[1][389] ;
  wire \shift_array_reg_n_0_[1][38] ;
  wire \shift_array_reg_n_0_[1][390] ;
  wire \shift_array_reg_n_0_[1][391] ;
  wire \shift_array_reg_n_0_[1][392] ;
  wire \shift_array_reg_n_0_[1][393] ;
  wire \shift_array_reg_n_0_[1][394] ;
  wire \shift_array_reg_n_0_[1][395] ;
  wire \shift_array_reg_n_0_[1][396] ;
  wire \shift_array_reg_n_0_[1][397] ;
  wire \shift_array_reg_n_0_[1][398] ;
  wire \shift_array_reg_n_0_[1][399] ;
  wire \shift_array_reg_n_0_[1][39] ;
  wire \shift_array_reg_n_0_[1][3] ;
  wire \shift_array_reg_n_0_[1][400] ;
  wire \shift_array_reg_n_0_[1][401] ;
  wire \shift_array_reg_n_0_[1][402] ;
  wire \shift_array_reg_n_0_[1][403] ;
  wire \shift_array_reg_n_0_[1][404] ;
  wire \shift_array_reg_n_0_[1][405] ;
  wire \shift_array_reg_n_0_[1][406] ;
  wire \shift_array_reg_n_0_[1][407] ;
  wire \shift_array_reg_n_0_[1][408] ;
  wire \shift_array_reg_n_0_[1][409] ;
  wire \shift_array_reg_n_0_[1][40] ;
  wire \shift_array_reg_n_0_[1][410] ;
  wire \shift_array_reg_n_0_[1][411] ;
  wire \shift_array_reg_n_0_[1][412] ;
  wire \shift_array_reg_n_0_[1][413] ;
  wire \shift_array_reg_n_0_[1][414] ;
  wire \shift_array_reg_n_0_[1][415] ;
  wire \shift_array_reg_n_0_[1][416] ;
  wire \shift_array_reg_n_0_[1][417] ;
  wire \shift_array_reg_n_0_[1][418] ;
  wire \shift_array_reg_n_0_[1][419] ;
  wire \shift_array_reg_n_0_[1][41] ;
  wire \shift_array_reg_n_0_[1][420] ;
  wire \shift_array_reg_n_0_[1][421] ;
  wire \shift_array_reg_n_0_[1][422] ;
  wire \shift_array_reg_n_0_[1][423] ;
  wire \shift_array_reg_n_0_[1][424] ;
  wire \shift_array_reg_n_0_[1][425] ;
  wire \shift_array_reg_n_0_[1][426] ;
  wire \shift_array_reg_n_0_[1][427] ;
  wire \shift_array_reg_n_0_[1][428] ;
  wire \shift_array_reg_n_0_[1][429] ;
  wire \shift_array_reg_n_0_[1][42] ;
  wire \shift_array_reg_n_0_[1][430] ;
  wire \shift_array_reg_n_0_[1][431] ;
  wire \shift_array_reg_n_0_[1][432] ;
  wire \shift_array_reg_n_0_[1][433] ;
  wire \shift_array_reg_n_0_[1][434] ;
  wire \shift_array_reg_n_0_[1][435] ;
  wire \shift_array_reg_n_0_[1][436] ;
  wire \shift_array_reg_n_0_[1][437] ;
  wire \shift_array_reg_n_0_[1][438] ;
  wire \shift_array_reg_n_0_[1][439] ;
  wire \shift_array_reg_n_0_[1][43] ;
  wire \shift_array_reg_n_0_[1][440] ;
  wire \shift_array_reg_n_0_[1][441] ;
  wire \shift_array_reg_n_0_[1][442] ;
  wire \shift_array_reg_n_0_[1][443] ;
  wire \shift_array_reg_n_0_[1][444] ;
  wire \shift_array_reg_n_0_[1][445] ;
  wire \shift_array_reg_n_0_[1][446] ;
  wire \shift_array_reg_n_0_[1][447] ;
  wire \shift_array_reg_n_0_[1][448] ;
  wire \shift_array_reg_n_0_[1][449] ;
  wire \shift_array_reg_n_0_[1][44] ;
  wire \shift_array_reg_n_0_[1][450] ;
  wire \shift_array_reg_n_0_[1][451] ;
  wire \shift_array_reg_n_0_[1][452] ;
  wire \shift_array_reg_n_0_[1][453] ;
  wire \shift_array_reg_n_0_[1][454] ;
  wire \shift_array_reg_n_0_[1][455] ;
  wire \shift_array_reg_n_0_[1][456] ;
  wire \shift_array_reg_n_0_[1][457] ;
  wire \shift_array_reg_n_0_[1][458] ;
  wire \shift_array_reg_n_0_[1][459] ;
  wire \shift_array_reg_n_0_[1][45] ;
  wire \shift_array_reg_n_0_[1][460] ;
  wire \shift_array_reg_n_0_[1][461] ;
  wire \shift_array_reg_n_0_[1][462] ;
  wire \shift_array_reg_n_0_[1][463] ;
  wire \shift_array_reg_n_0_[1][464] ;
  wire \shift_array_reg_n_0_[1][465] ;
  wire \shift_array_reg_n_0_[1][466] ;
  wire \shift_array_reg_n_0_[1][467] ;
  wire \shift_array_reg_n_0_[1][468] ;
  wire \shift_array_reg_n_0_[1][469] ;
  wire \shift_array_reg_n_0_[1][46] ;
  wire \shift_array_reg_n_0_[1][470] ;
  wire \shift_array_reg_n_0_[1][471] ;
  wire \shift_array_reg_n_0_[1][472] ;
  wire \shift_array_reg_n_0_[1][473] ;
  wire \shift_array_reg_n_0_[1][474] ;
  wire \shift_array_reg_n_0_[1][475] ;
  wire \shift_array_reg_n_0_[1][476] ;
  wire \shift_array_reg_n_0_[1][477] ;
  wire \shift_array_reg_n_0_[1][478] ;
  wire \shift_array_reg_n_0_[1][479] ;
  wire \shift_array_reg_n_0_[1][47] ;
  wire \shift_array_reg_n_0_[1][480] ;
  wire \shift_array_reg_n_0_[1][481] ;
  wire \shift_array_reg_n_0_[1][482] ;
  wire \shift_array_reg_n_0_[1][483] ;
  wire \shift_array_reg_n_0_[1][484] ;
  wire \shift_array_reg_n_0_[1][485] ;
  wire \shift_array_reg_n_0_[1][486] ;
  wire \shift_array_reg_n_0_[1][487] ;
  wire \shift_array_reg_n_0_[1][488] ;
  wire \shift_array_reg_n_0_[1][489] ;
  wire \shift_array_reg_n_0_[1][48] ;
  wire \shift_array_reg_n_0_[1][490] ;
  wire \shift_array_reg_n_0_[1][491] ;
  wire \shift_array_reg_n_0_[1][492] ;
  wire \shift_array_reg_n_0_[1][493] ;
  wire \shift_array_reg_n_0_[1][494] ;
  wire \shift_array_reg_n_0_[1][495] ;
  wire \shift_array_reg_n_0_[1][496] ;
  wire \shift_array_reg_n_0_[1][497] ;
  wire \shift_array_reg_n_0_[1][498] ;
  wire \shift_array_reg_n_0_[1][499] ;
  wire \shift_array_reg_n_0_[1][49] ;
  wire \shift_array_reg_n_0_[1][4] ;
  wire \shift_array_reg_n_0_[1][500] ;
  wire \shift_array_reg_n_0_[1][501] ;
  wire \shift_array_reg_n_0_[1][502] ;
  wire \shift_array_reg_n_0_[1][503] ;
  wire \shift_array_reg_n_0_[1][504] ;
  wire \shift_array_reg_n_0_[1][505] ;
  wire \shift_array_reg_n_0_[1][506] ;
  wire \shift_array_reg_n_0_[1][507] ;
  wire \shift_array_reg_n_0_[1][508] ;
  wire \shift_array_reg_n_0_[1][509] ;
  wire \shift_array_reg_n_0_[1][50] ;
  wire \shift_array_reg_n_0_[1][510] ;
  wire \shift_array_reg_n_0_[1][511] ;
  wire \shift_array_reg_n_0_[1][512] ;
  wire \shift_array_reg_n_0_[1][513] ;
  wire \shift_array_reg_n_0_[1][514] ;
  wire \shift_array_reg_n_0_[1][515] ;
  wire \shift_array_reg_n_0_[1][516] ;
  wire \shift_array_reg_n_0_[1][517] ;
  wire \shift_array_reg_n_0_[1][518] ;
  wire \shift_array_reg_n_0_[1][519] ;
  wire \shift_array_reg_n_0_[1][51] ;
  wire \shift_array_reg_n_0_[1][520] ;
  wire \shift_array_reg_n_0_[1][521] ;
  wire \shift_array_reg_n_0_[1][522] ;
  wire \shift_array_reg_n_0_[1][523] ;
  wire \shift_array_reg_n_0_[1][524] ;
  wire \shift_array_reg_n_0_[1][525] ;
  wire \shift_array_reg_n_0_[1][526] ;
  wire \shift_array_reg_n_0_[1][527] ;
  wire \shift_array_reg_n_0_[1][528] ;
  wire \shift_array_reg_n_0_[1][529] ;
  wire \shift_array_reg_n_0_[1][52] ;
  wire \shift_array_reg_n_0_[1][530] ;
  wire \shift_array_reg_n_0_[1][531] ;
  wire \shift_array_reg_n_0_[1][532] ;
  wire \shift_array_reg_n_0_[1][533] ;
  wire \shift_array_reg_n_0_[1][534] ;
  wire \shift_array_reg_n_0_[1][535] ;
  wire \shift_array_reg_n_0_[1][536] ;
  wire \shift_array_reg_n_0_[1][537] ;
  wire \shift_array_reg_n_0_[1][538] ;
  wire \shift_array_reg_n_0_[1][539] ;
  wire \shift_array_reg_n_0_[1][53] ;
  wire \shift_array_reg_n_0_[1][540] ;
  wire \shift_array_reg_n_0_[1][541] ;
  wire \shift_array_reg_n_0_[1][542] ;
  wire \shift_array_reg_n_0_[1][543] ;
  wire \shift_array_reg_n_0_[1][544] ;
  wire \shift_array_reg_n_0_[1][545] ;
  wire \shift_array_reg_n_0_[1][546] ;
  wire \shift_array_reg_n_0_[1][547] ;
  wire \shift_array_reg_n_0_[1][548] ;
  wire \shift_array_reg_n_0_[1][549] ;
  wire \shift_array_reg_n_0_[1][54] ;
  wire \shift_array_reg_n_0_[1][550] ;
  wire \shift_array_reg_n_0_[1][551] ;
  wire \shift_array_reg_n_0_[1][552] ;
  wire \shift_array_reg_n_0_[1][553] ;
  wire \shift_array_reg_n_0_[1][554] ;
  wire \shift_array_reg_n_0_[1][555] ;
  wire \shift_array_reg_n_0_[1][556] ;
  wire \shift_array_reg_n_0_[1][557] ;
  wire \shift_array_reg_n_0_[1][558] ;
  wire \shift_array_reg_n_0_[1][559] ;
  wire \shift_array_reg_n_0_[1][55] ;
  wire \shift_array_reg_n_0_[1][560] ;
  wire \shift_array_reg_n_0_[1][561] ;
  wire \shift_array_reg_n_0_[1][562] ;
  wire \shift_array_reg_n_0_[1][563] ;
  wire \shift_array_reg_n_0_[1][564] ;
  wire \shift_array_reg_n_0_[1][565] ;
  wire \shift_array_reg_n_0_[1][566] ;
  wire \shift_array_reg_n_0_[1][567] ;
  wire \shift_array_reg_n_0_[1][568] ;
  wire \shift_array_reg_n_0_[1][569] ;
  wire \shift_array_reg_n_0_[1][56] ;
  wire \shift_array_reg_n_0_[1][570] ;
  wire \shift_array_reg_n_0_[1][571] ;
  wire \shift_array_reg_n_0_[1][572] ;
  wire \shift_array_reg_n_0_[1][573] ;
  wire \shift_array_reg_n_0_[1][574] ;
  wire \shift_array_reg_n_0_[1][575] ;
  wire \shift_array_reg_n_0_[1][576] ;
  wire \shift_array_reg_n_0_[1][577] ;
  wire \shift_array_reg_n_0_[1][578] ;
  wire \shift_array_reg_n_0_[1][579] ;
  wire \shift_array_reg_n_0_[1][57] ;
  wire \shift_array_reg_n_0_[1][580] ;
  wire \shift_array_reg_n_0_[1][581] ;
  wire \shift_array_reg_n_0_[1][582] ;
  wire \shift_array_reg_n_0_[1][583] ;
  wire \shift_array_reg_n_0_[1][584] ;
  wire \shift_array_reg_n_0_[1][585] ;
  wire \shift_array_reg_n_0_[1][586] ;
  wire \shift_array_reg_n_0_[1][587] ;
  wire \shift_array_reg_n_0_[1][588] ;
  wire \shift_array_reg_n_0_[1][589] ;
  wire \shift_array_reg_n_0_[1][58] ;
  wire \shift_array_reg_n_0_[1][590] ;
  wire \shift_array_reg_n_0_[1][591] ;
  wire \shift_array_reg_n_0_[1][592] ;
  wire \shift_array_reg_n_0_[1][593] ;
  wire \shift_array_reg_n_0_[1][594] ;
  wire \shift_array_reg_n_0_[1][595] ;
  wire \shift_array_reg_n_0_[1][596] ;
  wire \shift_array_reg_n_0_[1][597] ;
  wire \shift_array_reg_n_0_[1][598] ;
  wire \shift_array_reg_n_0_[1][599] ;
  wire \shift_array_reg_n_0_[1][59] ;
  wire \shift_array_reg_n_0_[1][5] ;
  wire \shift_array_reg_n_0_[1][600] ;
  wire \shift_array_reg_n_0_[1][601] ;
  wire \shift_array_reg_n_0_[1][602] ;
  wire \shift_array_reg_n_0_[1][603] ;
  wire \shift_array_reg_n_0_[1][604] ;
  wire \shift_array_reg_n_0_[1][605] ;
  wire \shift_array_reg_n_0_[1][606] ;
  wire \shift_array_reg_n_0_[1][607] ;
  wire \shift_array_reg_n_0_[1][608] ;
  wire \shift_array_reg_n_0_[1][609] ;
  wire \shift_array_reg_n_0_[1][60] ;
  wire \shift_array_reg_n_0_[1][610] ;
  wire \shift_array_reg_n_0_[1][611] ;
  wire \shift_array_reg_n_0_[1][612] ;
  wire \shift_array_reg_n_0_[1][613] ;
  wire \shift_array_reg_n_0_[1][614] ;
  wire \shift_array_reg_n_0_[1][615] ;
  wire \shift_array_reg_n_0_[1][616] ;
  wire \shift_array_reg_n_0_[1][617] ;
  wire \shift_array_reg_n_0_[1][618] ;
  wire \shift_array_reg_n_0_[1][619] ;
  wire \shift_array_reg_n_0_[1][61] ;
  wire \shift_array_reg_n_0_[1][620] ;
  wire \shift_array_reg_n_0_[1][621] ;
  wire \shift_array_reg_n_0_[1][622] ;
  wire \shift_array_reg_n_0_[1][623] ;
  wire \shift_array_reg_n_0_[1][624] ;
  wire \shift_array_reg_n_0_[1][625] ;
  wire \shift_array_reg_n_0_[1][626] ;
  wire \shift_array_reg_n_0_[1][627] ;
  wire \shift_array_reg_n_0_[1][628] ;
  wire \shift_array_reg_n_0_[1][629] ;
  wire \shift_array_reg_n_0_[1][62] ;
  wire \shift_array_reg_n_0_[1][630] ;
  wire \shift_array_reg_n_0_[1][631] ;
  wire \shift_array_reg_n_0_[1][632] ;
  wire \shift_array_reg_n_0_[1][633] ;
  wire \shift_array_reg_n_0_[1][634] ;
  wire \shift_array_reg_n_0_[1][635] ;
  wire \shift_array_reg_n_0_[1][636] ;
  wire \shift_array_reg_n_0_[1][637] ;
  wire \shift_array_reg_n_0_[1][638] ;
  wire \shift_array_reg_n_0_[1][639] ;
  wire \shift_array_reg_n_0_[1][63] ;
  wire \shift_array_reg_n_0_[1][640] ;
  wire \shift_array_reg_n_0_[1][641] ;
  wire \shift_array_reg_n_0_[1][642] ;
  wire \shift_array_reg_n_0_[1][643] ;
  wire \shift_array_reg_n_0_[1][644] ;
  wire \shift_array_reg_n_0_[1][645] ;
  wire \shift_array_reg_n_0_[1][646] ;
  wire \shift_array_reg_n_0_[1][647] ;
  wire \shift_array_reg_n_0_[1][648] ;
  wire \shift_array_reg_n_0_[1][649] ;
  wire \shift_array_reg_n_0_[1][64] ;
  wire \shift_array_reg_n_0_[1][650] ;
  wire \shift_array_reg_n_0_[1][651] ;
  wire \shift_array_reg_n_0_[1][652] ;
  wire \shift_array_reg_n_0_[1][653] ;
  wire \shift_array_reg_n_0_[1][654] ;
  wire \shift_array_reg_n_0_[1][655] ;
  wire \shift_array_reg_n_0_[1][656] ;
  wire \shift_array_reg_n_0_[1][657] ;
  wire \shift_array_reg_n_0_[1][658] ;
  wire \shift_array_reg_n_0_[1][659] ;
  wire \shift_array_reg_n_0_[1][65] ;
  wire \shift_array_reg_n_0_[1][660] ;
  wire \shift_array_reg_n_0_[1][661] ;
  wire \shift_array_reg_n_0_[1][662] ;
  wire \shift_array_reg_n_0_[1][663] ;
  wire \shift_array_reg_n_0_[1][664] ;
  wire \shift_array_reg_n_0_[1][665] ;
  wire \shift_array_reg_n_0_[1][666] ;
  wire \shift_array_reg_n_0_[1][667] ;
  wire \shift_array_reg_n_0_[1][668] ;
  wire \shift_array_reg_n_0_[1][669] ;
  wire \shift_array_reg_n_0_[1][66] ;
  wire \shift_array_reg_n_0_[1][670] ;
  wire \shift_array_reg_n_0_[1][671] ;
  wire \shift_array_reg_n_0_[1][672] ;
  wire \shift_array_reg_n_0_[1][673] ;
  wire \shift_array_reg_n_0_[1][674] ;
  wire \shift_array_reg_n_0_[1][675] ;
  wire \shift_array_reg_n_0_[1][676] ;
  wire \shift_array_reg_n_0_[1][677] ;
  wire \shift_array_reg_n_0_[1][678] ;
  wire \shift_array_reg_n_0_[1][679] ;
  wire \shift_array_reg_n_0_[1][67] ;
  wire \shift_array_reg_n_0_[1][680] ;
  wire \shift_array_reg_n_0_[1][681] ;
  wire \shift_array_reg_n_0_[1][682] ;
  wire \shift_array_reg_n_0_[1][683] ;
  wire \shift_array_reg_n_0_[1][684] ;
  wire \shift_array_reg_n_0_[1][685] ;
  wire \shift_array_reg_n_0_[1][686] ;
  wire \shift_array_reg_n_0_[1][687] ;
  wire \shift_array_reg_n_0_[1][688] ;
  wire \shift_array_reg_n_0_[1][689] ;
  wire \shift_array_reg_n_0_[1][68] ;
  wire \shift_array_reg_n_0_[1][690] ;
  wire \shift_array_reg_n_0_[1][691] ;
  wire \shift_array_reg_n_0_[1][692] ;
  wire \shift_array_reg_n_0_[1][693] ;
  wire \shift_array_reg_n_0_[1][694] ;
  wire \shift_array_reg_n_0_[1][695] ;
  wire \shift_array_reg_n_0_[1][696] ;
  wire \shift_array_reg_n_0_[1][697] ;
  wire \shift_array_reg_n_0_[1][698] ;
  wire \shift_array_reg_n_0_[1][699] ;
  wire \shift_array_reg_n_0_[1][69] ;
  wire \shift_array_reg_n_0_[1][6] ;
  wire \shift_array_reg_n_0_[1][700] ;
  wire \shift_array_reg_n_0_[1][701] ;
  wire \shift_array_reg_n_0_[1][702] ;
  wire \shift_array_reg_n_0_[1][703] ;
  wire \shift_array_reg_n_0_[1][704] ;
  wire \shift_array_reg_n_0_[1][705] ;
  wire \shift_array_reg_n_0_[1][706] ;
  wire \shift_array_reg_n_0_[1][707] ;
  wire \shift_array_reg_n_0_[1][708] ;
  wire \shift_array_reg_n_0_[1][709] ;
  wire \shift_array_reg_n_0_[1][70] ;
  wire \shift_array_reg_n_0_[1][710] ;
  wire \shift_array_reg_n_0_[1][711] ;
  wire \shift_array_reg_n_0_[1][712] ;
  wire \shift_array_reg_n_0_[1][713] ;
  wire \shift_array_reg_n_0_[1][714] ;
  wire \shift_array_reg_n_0_[1][715] ;
  wire \shift_array_reg_n_0_[1][716] ;
  wire \shift_array_reg_n_0_[1][717] ;
  wire \shift_array_reg_n_0_[1][718] ;
  wire \shift_array_reg_n_0_[1][719] ;
  wire \shift_array_reg_n_0_[1][71] ;
  wire \shift_array_reg_n_0_[1][720] ;
  wire \shift_array_reg_n_0_[1][721] ;
  wire \shift_array_reg_n_0_[1][722] ;
  wire \shift_array_reg_n_0_[1][723] ;
  wire \shift_array_reg_n_0_[1][724] ;
  wire \shift_array_reg_n_0_[1][725] ;
  wire \shift_array_reg_n_0_[1][726] ;
  wire \shift_array_reg_n_0_[1][727] ;
  wire \shift_array_reg_n_0_[1][728] ;
  wire \shift_array_reg_n_0_[1][729] ;
  wire \shift_array_reg_n_0_[1][72] ;
  wire \shift_array_reg_n_0_[1][730] ;
  wire \shift_array_reg_n_0_[1][731] ;
  wire \shift_array_reg_n_0_[1][732] ;
  wire \shift_array_reg_n_0_[1][733] ;
  wire \shift_array_reg_n_0_[1][734] ;
  wire \shift_array_reg_n_0_[1][735] ;
  wire \shift_array_reg_n_0_[1][736] ;
  wire \shift_array_reg_n_0_[1][737] ;
  wire \shift_array_reg_n_0_[1][738] ;
  wire \shift_array_reg_n_0_[1][739] ;
  wire \shift_array_reg_n_0_[1][73] ;
  wire \shift_array_reg_n_0_[1][740] ;
  wire \shift_array_reg_n_0_[1][741] ;
  wire \shift_array_reg_n_0_[1][742] ;
  wire \shift_array_reg_n_0_[1][743] ;
  wire \shift_array_reg_n_0_[1][744] ;
  wire \shift_array_reg_n_0_[1][745] ;
  wire \shift_array_reg_n_0_[1][746] ;
  wire \shift_array_reg_n_0_[1][747] ;
  wire \shift_array_reg_n_0_[1][748] ;
  wire \shift_array_reg_n_0_[1][749] ;
  wire \shift_array_reg_n_0_[1][74] ;
  wire \shift_array_reg_n_0_[1][750] ;
  wire \shift_array_reg_n_0_[1][751] ;
  wire \shift_array_reg_n_0_[1][752] ;
  wire \shift_array_reg_n_0_[1][753] ;
  wire \shift_array_reg_n_0_[1][754] ;
  wire \shift_array_reg_n_0_[1][755] ;
  wire \shift_array_reg_n_0_[1][756] ;
  wire \shift_array_reg_n_0_[1][757] ;
  wire \shift_array_reg_n_0_[1][758] ;
  wire \shift_array_reg_n_0_[1][759] ;
  wire \shift_array_reg_n_0_[1][75] ;
  wire \shift_array_reg_n_0_[1][760] ;
  wire \shift_array_reg_n_0_[1][761] ;
  wire \shift_array_reg_n_0_[1][762] ;
  wire \shift_array_reg_n_0_[1][763] ;
  wire \shift_array_reg_n_0_[1][764] ;
  wire \shift_array_reg_n_0_[1][765] ;
  wire \shift_array_reg_n_0_[1][766] ;
  wire \shift_array_reg_n_0_[1][767] ;
  wire \shift_array_reg_n_0_[1][768] ;
  wire \shift_array_reg_n_0_[1][769] ;
  wire \shift_array_reg_n_0_[1][76] ;
  wire \shift_array_reg_n_0_[1][770] ;
  wire \shift_array_reg_n_0_[1][771] ;
  wire \shift_array_reg_n_0_[1][772] ;
  wire \shift_array_reg_n_0_[1][773] ;
  wire \shift_array_reg_n_0_[1][774] ;
  wire \shift_array_reg_n_0_[1][775] ;
  wire \shift_array_reg_n_0_[1][776] ;
  wire \shift_array_reg_n_0_[1][777] ;
  wire \shift_array_reg_n_0_[1][778] ;
  wire \shift_array_reg_n_0_[1][779] ;
  wire \shift_array_reg_n_0_[1][77] ;
  wire \shift_array_reg_n_0_[1][780] ;
  wire \shift_array_reg_n_0_[1][781] ;
  wire \shift_array_reg_n_0_[1][782] ;
  wire \shift_array_reg_n_0_[1][783] ;
  wire \shift_array_reg_n_0_[1][784] ;
  wire \shift_array_reg_n_0_[1][785] ;
  wire \shift_array_reg_n_0_[1][786] ;
  wire \shift_array_reg_n_0_[1][787] ;
  wire \shift_array_reg_n_0_[1][788] ;
  wire \shift_array_reg_n_0_[1][789] ;
  wire \shift_array_reg_n_0_[1][78] ;
  wire \shift_array_reg_n_0_[1][790] ;
  wire \shift_array_reg_n_0_[1][791] ;
  wire \shift_array_reg_n_0_[1][792] ;
  wire \shift_array_reg_n_0_[1][793] ;
  wire \shift_array_reg_n_0_[1][794] ;
  wire \shift_array_reg_n_0_[1][795] ;
  wire \shift_array_reg_n_0_[1][796] ;
  wire \shift_array_reg_n_0_[1][797] ;
  wire \shift_array_reg_n_0_[1][798] ;
  wire \shift_array_reg_n_0_[1][799] ;
  wire \shift_array_reg_n_0_[1][79] ;
  wire \shift_array_reg_n_0_[1][7] ;
  wire \shift_array_reg_n_0_[1][800] ;
  wire \shift_array_reg_n_0_[1][801] ;
  wire \shift_array_reg_n_0_[1][802] ;
  wire \shift_array_reg_n_0_[1][803] ;
  wire \shift_array_reg_n_0_[1][804] ;
  wire \shift_array_reg_n_0_[1][805] ;
  wire \shift_array_reg_n_0_[1][806] ;
  wire \shift_array_reg_n_0_[1][807] ;
  wire \shift_array_reg_n_0_[1][808] ;
  wire \shift_array_reg_n_0_[1][809] ;
  wire \shift_array_reg_n_0_[1][80] ;
  wire \shift_array_reg_n_0_[1][810] ;
  wire \shift_array_reg_n_0_[1][811] ;
  wire \shift_array_reg_n_0_[1][812] ;
  wire \shift_array_reg_n_0_[1][813] ;
  wire \shift_array_reg_n_0_[1][814] ;
  wire \shift_array_reg_n_0_[1][815] ;
  wire \shift_array_reg_n_0_[1][816] ;
  wire \shift_array_reg_n_0_[1][817] ;
  wire \shift_array_reg_n_0_[1][818] ;
  wire \shift_array_reg_n_0_[1][819] ;
  wire \shift_array_reg_n_0_[1][81] ;
  wire \shift_array_reg_n_0_[1][820] ;
  wire \shift_array_reg_n_0_[1][821] ;
  wire \shift_array_reg_n_0_[1][822] ;
  wire \shift_array_reg_n_0_[1][823] ;
  wire \shift_array_reg_n_0_[1][824] ;
  wire \shift_array_reg_n_0_[1][825] ;
  wire \shift_array_reg_n_0_[1][826] ;
  wire \shift_array_reg_n_0_[1][827] ;
  wire \shift_array_reg_n_0_[1][828] ;
  wire \shift_array_reg_n_0_[1][829] ;
  wire \shift_array_reg_n_0_[1][82] ;
  wire \shift_array_reg_n_0_[1][830] ;
  wire \shift_array_reg_n_0_[1][831] ;
  wire \shift_array_reg_n_0_[1][832] ;
  wire \shift_array_reg_n_0_[1][833] ;
  wire \shift_array_reg_n_0_[1][834] ;
  wire \shift_array_reg_n_0_[1][835] ;
  wire \shift_array_reg_n_0_[1][836] ;
  wire \shift_array_reg_n_0_[1][837] ;
  wire \shift_array_reg_n_0_[1][838] ;
  wire \shift_array_reg_n_0_[1][839] ;
  wire \shift_array_reg_n_0_[1][83] ;
  wire \shift_array_reg_n_0_[1][840] ;
  wire \shift_array_reg_n_0_[1][841] ;
  wire \shift_array_reg_n_0_[1][842] ;
  wire \shift_array_reg_n_0_[1][843] ;
  wire \shift_array_reg_n_0_[1][844] ;
  wire \shift_array_reg_n_0_[1][845] ;
  wire \shift_array_reg_n_0_[1][846] ;
  wire \shift_array_reg_n_0_[1][847] ;
  wire \shift_array_reg_n_0_[1][848] ;
  wire \shift_array_reg_n_0_[1][849] ;
  wire \shift_array_reg_n_0_[1][84] ;
  wire \shift_array_reg_n_0_[1][850] ;
  wire \shift_array_reg_n_0_[1][851] ;
  wire \shift_array_reg_n_0_[1][852] ;
  wire \shift_array_reg_n_0_[1][853] ;
  wire \shift_array_reg_n_0_[1][854] ;
  wire \shift_array_reg_n_0_[1][855] ;
  wire \shift_array_reg_n_0_[1][856] ;
  wire \shift_array_reg_n_0_[1][857] ;
  wire \shift_array_reg_n_0_[1][858] ;
  wire \shift_array_reg_n_0_[1][859] ;
  wire \shift_array_reg_n_0_[1][85] ;
  wire \shift_array_reg_n_0_[1][860] ;
  wire \shift_array_reg_n_0_[1][861] ;
  wire \shift_array_reg_n_0_[1][862] ;
  wire \shift_array_reg_n_0_[1][863] ;
  wire \shift_array_reg_n_0_[1][864] ;
  wire \shift_array_reg_n_0_[1][865] ;
  wire \shift_array_reg_n_0_[1][866] ;
  wire \shift_array_reg_n_0_[1][867] ;
  wire \shift_array_reg_n_0_[1][868] ;
  wire \shift_array_reg_n_0_[1][869] ;
  wire \shift_array_reg_n_0_[1][86] ;
  wire \shift_array_reg_n_0_[1][870] ;
  wire \shift_array_reg_n_0_[1][871] ;
  wire \shift_array_reg_n_0_[1][872] ;
  wire \shift_array_reg_n_0_[1][873] ;
  wire \shift_array_reg_n_0_[1][874] ;
  wire \shift_array_reg_n_0_[1][875] ;
  wire \shift_array_reg_n_0_[1][876] ;
  wire \shift_array_reg_n_0_[1][877] ;
  wire \shift_array_reg_n_0_[1][878] ;
  wire \shift_array_reg_n_0_[1][879] ;
  wire \shift_array_reg_n_0_[1][87] ;
  wire \shift_array_reg_n_0_[1][880] ;
  wire \shift_array_reg_n_0_[1][881] ;
  wire \shift_array_reg_n_0_[1][882] ;
  wire \shift_array_reg_n_0_[1][883] ;
  wire \shift_array_reg_n_0_[1][884] ;
  wire \shift_array_reg_n_0_[1][885] ;
  wire \shift_array_reg_n_0_[1][886] ;
  wire \shift_array_reg_n_0_[1][887] ;
  wire \shift_array_reg_n_0_[1][888] ;
  wire \shift_array_reg_n_0_[1][889] ;
  wire \shift_array_reg_n_0_[1][88] ;
  wire \shift_array_reg_n_0_[1][890] ;
  wire \shift_array_reg_n_0_[1][891] ;
  wire \shift_array_reg_n_0_[1][892] ;
  wire \shift_array_reg_n_0_[1][893] ;
  wire \shift_array_reg_n_0_[1][894] ;
  wire \shift_array_reg_n_0_[1][895] ;
  wire \shift_array_reg_n_0_[1][896] ;
  wire \shift_array_reg_n_0_[1][897] ;
  wire \shift_array_reg_n_0_[1][898] ;
  wire \shift_array_reg_n_0_[1][899] ;
  wire \shift_array_reg_n_0_[1][89] ;
  wire \shift_array_reg_n_0_[1][8] ;
  wire \shift_array_reg_n_0_[1][900] ;
  wire \shift_array_reg_n_0_[1][901] ;
  wire \shift_array_reg_n_0_[1][902] ;
  wire \shift_array_reg_n_0_[1][903] ;
  wire \shift_array_reg_n_0_[1][904] ;
  wire \shift_array_reg_n_0_[1][905] ;
  wire \shift_array_reg_n_0_[1][906] ;
  wire \shift_array_reg_n_0_[1][907] ;
  wire \shift_array_reg_n_0_[1][908] ;
  wire \shift_array_reg_n_0_[1][909] ;
  wire \shift_array_reg_n_0_[1][90] ;
  wire \shift_array_reg_n_0_[1][910] ;
  wire \shift_array_reg_n_0_[1][911] ;
  wire \shift_array_reg_n_0_[1][912] ;
  wire \shift_array_reg_n_0_[1][913] ;
  wire \shift_array_reg_n_0_[1][914] ;
  wire \shift_array_reg_n_0_[1][915] ;
  wire \shift_array_reg_n_0_[1][916] ;
  wire \shift_array_reg_n_0_[1][917] ;
  wire \shift_array_reg_n_0_[1][918] ;
  wire \shift_array_reg_n_0_[1][919] ;
  wire \shift_array_reg_n_0_[1][91] ;
  wire \shift_array_reg_n_0_[1][920] ;
  wire \shift_array_reg_n_0_[1][921] ;
  wire \shift_array_reg_n_0_[1][922] ;
  wire \shift_array_reg_n_0_[1][923] ;
  wire \shift_array_reg_n_0_[1][924] ;
  wire \shift_array_reg_n_0_[1][925] ;
  wire \shift_array_reg_n_0_[1][926] ;
  wire \shift_array_reg_n_0_[1][927] ;
  wire \shift_array_reg_n_0_[1][928] ;
  wire \shift_array_reg_n_0_[1][929] ;
  wire \shift_array_reg_n_0_[1][92] ;
  wire \shift_array_reg_n_0_[1][930] ;
  wire \shift_array_reg_n_0_[1][931] ;
  wire \shift_array_reg_n_0_[1][932] ;
  wire \shift_array_reg_n_0_[1][933] ;
  wire \shift_array_reg_n_0_[1][934] ;
  wire \shift_array_reg_n_0_[1][935] ;
  wire \shift_array_reg_n_0_[1][936] ;
  wire \shift_array_reg_n_0_[1][937] ;
  wire \shift_array_reg_n_0_[1][938] ;
  wire \shift_array_reg_n_0_[1][939] ;
  wire \shift_array_reg_n_0_[1][93] ;
  wire \shift_array_reg_n_0_[1][940] ;
  wire \shift_array_reg_n_0_[1][941] ;
  wire \shift_array_reg_n_0_[1][942] ;
  wire \shift_array_reg_n_0_[1][943] ;
  wire \shift_array_reg_n_0_[1][944] ;
  wire \shift_array_reg_n_0_[1][945] ;
  wire \shift_array_reg_n_0_[1][946] ;
  wire \shift_array_reg_n_0_[1][947] ;
  wire \shift_array_reg_n_0_[1][948] ;
  wire \shift_array_reg_n_0_[1][949] ;
  wire \shift_array_reg_n_0_[1][94] ;
  wire \shift_array_reg_n_0_[1][950] ;
  wire \shift_array_reg_n_0_[1][951] ;
  wire \shift_array_reg_n_0_[1][952] ;
  wire \shift_array_reg_n_0_[1][953] ;
  wire \shift_array_reg_n_0_[1][954] ;
  wire \shift_array_reg_n_0_[1][955] ;
  wire \shift_array_reg_n_0_[1][956] ;
  wire \shift_array_reg_n_0_[1][957] ;
  wire \shift_array_reg_n_0_[1][958] ;
  wire \shift_array_reg_n_0_[1][959] ;
  wire \shift_array_reg_n_0_[1][95] ;
  wire \shift_array_reg_n_0_[1][960] ;
  wire \shift_array_reg_n_0_[1][961] ;
  wire \shift_array_reg_n_0_[1][962] ;
  wire \shift_array_reg_n_0_[1][963] ;
  wire \shift_array_reg_n_0_[1][964] ;
  wire \shift_array_reg_n_0_[1][965] ;
  wire \shift_array_reg_n_0_[1][966] ;
  wire \shift_array_reg_n_0_[1][967] ;
  wire \shift_array_reg_n_0_[1][968] ;
  wire \shift_array_reg_n_0_[1][969] ;
  wire \shift_array_reg_n_0_[1][96] ;
  wire \shift_array_reg_n_0_[1][970] ;
  wire \shift_array_reg_n_0_[1][971] ;
  wire \shift_array_reg_n_0_[1][972] ;
  wire \shift_array_reg_n_0_[1][973] ;
  wire \shift_array_reg_n_0_[1][974] ;
  wire \shift_array_reg_n_0_[1][975] ;
  wire \shift_array_reg_n_0_[1][976] ;
  wire \shift_array_reg_n_0_[1][977] ;
  wire \shift_array_reg_n_0_[1][978] ;
  wire \shift_array_reg_n_0_[1][979] ;
  wire \shift_array_reg_n_0_[1][97] ;
  wire \shift_array_reg_n_0_[1][980] ;
  wire \shift_array_reg_n_0_[1][981] ;
  wire \shift_array_reg_n_0_[1][982] ;
  wire \shift_array_reg_n_0_[1][983] ;
  wire \shift_array_reg_n_0_[1][984] ;
  wire \shift_array_reg_n_0_[1][985] ;
  wire \shift_array_reg_n_0_[1][986] ;
  wire \shift_array_reg_n_0_[1][987] ;
  wire \shift_array_reg_n_0_[1][988] ;
  wire \shift_array_reg_n_0_[1][989] ;
  wire \shift_array_reg_n_0_[1][98] ;
  wire \shift_array_reg_n_0_[1][990] ;
  wire \shift_array_reg_n_0_[1][991] ;
  wire \shift_array_reg_n_0_[1][992] ;
  wire \shift_array_reg_n_0_[1][993] ;
  wire \shift_array_reg_n_0_[1][994] ;
  wire \shift_array_reg_n_0_[1][995] ;
  wire \shift_array_reg_n_0_[1][996] ;
  wire \shift_array_reg_n_0_[1][997] ;
  wire \shift_array_reg_n_0_[1][998] ;
  wire \shift_array_reg_n_0_[1][999] ;
  wire \shift_array_reg_n_0_[1][99] ;
  wire \shift_array_reg_n_0_[1][9] ;

  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][0]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][0]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][0] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][0]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1000]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1000]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1000] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1000]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1001]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1001]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1001] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1001]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1002]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1002]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1002] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1002]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1003]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1003]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1003] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1003]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1004]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1004]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1004] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1004]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1005]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1005]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1005] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1005]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1006]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1006]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1006] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1006]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1007]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1007]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1007] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1007]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1008]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1008]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1008] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1008]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1009]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1009]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1009] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1009]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][100]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][100]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][100] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][100]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1010]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1010]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1010] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1010]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1011]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1011]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1011] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1011]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1012]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1012]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1012] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1012]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1013]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1013]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1013] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1013]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1014]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1014]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1014] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1014]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1015]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1015]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1015] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1015]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1016]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1016]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1016] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1016]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1017]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1017]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1017] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1017]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1018]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1018]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1018] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1018]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1019]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1019]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1019] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1019]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][101]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][101]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][101] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][101]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1020]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1020]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1020] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1020]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1021]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1021]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1021] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1021]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1022]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1022]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1022] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1022]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1023]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1023]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1023] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1023]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1024]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1024]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1024] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1024]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1025]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1025]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1025] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1025]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1026]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1026]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1026] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1026]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1027]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1027]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1027] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1027]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1028]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1028]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1028] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1028]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1029]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1029]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1029] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1029]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][102]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][102]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][102] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][102]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1030]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1030]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1030] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1030]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1031]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1031]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1031] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1031]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1032]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1032]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1032] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1032]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1033]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1033]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1033] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1033]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1034]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1034]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1034] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1034]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1035]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1035]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1035] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1035]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1036]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1036]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1036] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1036]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1037]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1037]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1037] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1037]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1038]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1038]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1038] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1038]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1039]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1039]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1039] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1039]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][103]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][103]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][103] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][103]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1040]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1040]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1040] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1040]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1041]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1041]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1041] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1041]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1042]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1042]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1042] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1042]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1043]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1043]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1043] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1043]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1044]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1044]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1044] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1044]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1045]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1045]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1045] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1045]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1046]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1046]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1046] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1046]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1047]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1047]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1047] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1047]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1048]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1048]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1048] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1048]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1049]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1049]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1049] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1049]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][104]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][104]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][104] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][104]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1050]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1050]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1050] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1050]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1051]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1051]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1051] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1051]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1052]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1052]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1052] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1052]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1053]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1053]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1053] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1053]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1054]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1054]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1054] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1054]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1055]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1055]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1055] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1055]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1056]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1056]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1056] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1056]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1057]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1057]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1057] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1057]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1058]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1058]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1058] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1058]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1059]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1059]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1059] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1059]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][105]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][105]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][105] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][105]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1060]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1060]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1060] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1060]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1061]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1061]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1061] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1061]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1062]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1062]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1062] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1062]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1063]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1063]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1063] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1063]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1064]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1064]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1064] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1064]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1065]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1065]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1065] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1065]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1066]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1066]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1066] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1066]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1067]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1067]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1067] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1067]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1068]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1068]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1068] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1068]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1069]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1069]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1069] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1069]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][106]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][106]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][106] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][106]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1070]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1070]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1070] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1070]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1071]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1071]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1071] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1071]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1072]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1072]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1072] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1072]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1073]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1073]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1073] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1073]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1074]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1074]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1074] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1074]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1075]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1075]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1075] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1075]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1076]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1076]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1076] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1076]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1077]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1077]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1077] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1077]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1078]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1078]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1078] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1078]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1079]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1079]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1079] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1079]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][107]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][107]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][107] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][107]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1080]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1080]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1080] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1080]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1081]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1081]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1081] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1081]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1082]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1082]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1082] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1082]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1083]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1083]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1083] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1083]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1084]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1084]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1084] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1084]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1085]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1085]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1085] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1085]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1086]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1086]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1086] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1086]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1087]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1087]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1087] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1087]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1088]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1088]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1088] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1088]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1089]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1089]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1089] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1089]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][108]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][108]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][108] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][108]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1090]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1090]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1090] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1090]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1091]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1091]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1091] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1091]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1092]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1092]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1092] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1092]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1093]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1093]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1093] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1093]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1094]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1094]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1094] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1094]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1095]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1095]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1095] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1095]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1096]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1096]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1096] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1096]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1097]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1097]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1097] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1097]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1098]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1098]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1098] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1098]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1099]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1099]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1099] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1099]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][109]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][109]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][109] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][109]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][10]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][10]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][10] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][10]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1100]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1100]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1100] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1100]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1101]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1101]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1101] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1101]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1102]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1102]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1102] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1102]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1103]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1103]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1103] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1103]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1104]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1104]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1104] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1104]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1105]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1105]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1105] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1105]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1106]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1106]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1106] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1106]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1107]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1107]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1107] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1107]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1108]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1108]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1108] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1108]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1109]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1109]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1109] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1109]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][110]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][110]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][110] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][110]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1110]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1110]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1110] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1110]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1111]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1111]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1111] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1111]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1112]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1112]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1112] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1112]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1113]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1113]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1113] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1113]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1114]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1114]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1114] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1114]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1115]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1115]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1115] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1115]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1116]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1116]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1116] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1116]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1117]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1117]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1117] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1117]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1118]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1118]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1118] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1118]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1119]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1119]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1119] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1119]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][111]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][111]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][111] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][111]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1120]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1120]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1120] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1120]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1121]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1121]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1121] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1121]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1122]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1122]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1122] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1122]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1123]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1123]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1123] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1123]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1124]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1124]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1124] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1124]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1125]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1125]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1125] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1125]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1126]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1126]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1126] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1126]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1127]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1127]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1127] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1127]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1128]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1128]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1128] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1128]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1129]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1129]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1129] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1129]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][112]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][112]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][112] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][112]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1130]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1130]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1130] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1130]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1131]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1131]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1131] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1131]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1132]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1132]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1132] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1132]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1133]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1133]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1133] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1133]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1134]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1134]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1134] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1134]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1135]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1135]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1135] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1135]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1136]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1136]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1136] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1136]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1137]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1137]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1137] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1137]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1138]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1138]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1138] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1138]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1139]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1139]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1139] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1139]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][113]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][113]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][113] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][113]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1140]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1140]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1140] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1140]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1141]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1141]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1141] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1141]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1142]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1142]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1142] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1142]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1143]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1143]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1143] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1143]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1144]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1144]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1144] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1144]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1145]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1145]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1145] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1145]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1146]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1146]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1146] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1146]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1147]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1147]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1147] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1147]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1148]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1148]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1148] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1148]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1149]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1149]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1149] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1149]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][114]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][114]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][114] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][114]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1150]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1150]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1150] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1150]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1151]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1151]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1151] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1151]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1152]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1152]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1152] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1152]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1153]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1153]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1153] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1153]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1154]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1154]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1154] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1154]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1155]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1155]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1155] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1155]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1156]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1156]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1156] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1156]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1157]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1157]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1157] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1157]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1158]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1158]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1158] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1158]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1159]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1159]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1159] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1159]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][115]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][115]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][115] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][115]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1160]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1160]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1160] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1160]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1161]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1161]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1161] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1161]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1162]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1162]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1162] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1162]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1163]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1163]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1163] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1163]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][116]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][116]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][116] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][116]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][117]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][117]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][117] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][117]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][118]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][118]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][118] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][118]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][119]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][119]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][119] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][119]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][11]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][11]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][11] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][11]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][120]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][120]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][120] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][120]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][121]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][121]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][121] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][121]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][122]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][122]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][122] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][122]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][123]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][123]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][123] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][123]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][124]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][124]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][124] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][124]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][125]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][125]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][125] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][125]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][126]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][126]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][126] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][126]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][127]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][127]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][127] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][127]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][128]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][128]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][128] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][128]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][129]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][129]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][129] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][129]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][12]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][12]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][12] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][12]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][130]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][130]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][130] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][130]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][131]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][131]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][131] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][131]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][132]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][132]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][132] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][132]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][133]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][133]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][133] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][133]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][134]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][134]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][134] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][134]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][135]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][135]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][135] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][135]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][136]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][136]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][136] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][136]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][137]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][137]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][137] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][137]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][138]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][138]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][138] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][138]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][139]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][139]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][139] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][139]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][13]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][13]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][13] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][13]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][140]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][140]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][140] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][140]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][141]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][141]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][141] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][141]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][142]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][142]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][142] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][142]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][143]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][143]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][143] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][143]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][144]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][144]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][144] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][144]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][145]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][145]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][145] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][145]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][146]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][146]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][146] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][146]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][147]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][147]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][147] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][147]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][148]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][148]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][148] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][148]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][149]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][149]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][149] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][149]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][14]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][14]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][14] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][14]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][150]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][150]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][150] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][150]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][151]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][151]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][151] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][151]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][152]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][152]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][152] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][152]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][153]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][153]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][153] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][153]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][154]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][154]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][154] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][154]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][155]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][155]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][155] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][155]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][156]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][156]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][156] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][156]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][157]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][157]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][157] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][157]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][158]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][158]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][158] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][158]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][159]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][159]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][159] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][159]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][15]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][15]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][15] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][15]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][160]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][160]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][160] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][160]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][161]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][161]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][161] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][161]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][162]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][162]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][162] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][162]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][163]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][163]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][163] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][163]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][164]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][164]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][164] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][164]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][165]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][165]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][165] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][165]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][166]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][166]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][166] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][166]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][167]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][167]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][167] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][167]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][168]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][168]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][168] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][168]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][169]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][169]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][169] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][169]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][16]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][16]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][16] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][16]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][170]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][170]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][170] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][170]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][171]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][171]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][171] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][171]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][172]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][172]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][172] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][172]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][173]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][173]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][173] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][173]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][174]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][174]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][174] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][174]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][175]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][175]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][175] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][175]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][176]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][176]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][176] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][176]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][177]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][177]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][177] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][177]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][178]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][178]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][178] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][178]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][179]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][179]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][179] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][179]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][17]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][17]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][17] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][17]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][180]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][180]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][180] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][180]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][181]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][181]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][181] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][181]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][182]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][182]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][182] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][182]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][183]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][183]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][183] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][183]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][184]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][184]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][184] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][184]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][185]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][185]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][185] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][185]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][186]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][186]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][186] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][186]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][187]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][187]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][187] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][187]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][188]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][188]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][188] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][188]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][189]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][189]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][189] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][189]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][18]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][18]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][18] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][18]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][190]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][190]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][190] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][190]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][191]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][191]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][191] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][191]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][192]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][192]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][192] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][192]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][193]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][193]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][193] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][193]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][194]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][194]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][194] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][194]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][195]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][195]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][195] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][195]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][196]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][196]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][196] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][196]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][197]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][197]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][197] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][197]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][198]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][198]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][198] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][198]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][199]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][199]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][199] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][199]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][19]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][19]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][19] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][19]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][1]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][1]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][1] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][1]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][200]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][200]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][200] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][200]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][201]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][201]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][201] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][201]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][202]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][202]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][202] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][202]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][203]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][203]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][203] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][203]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][204]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][204]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][204] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][204]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][205]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][205]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][205] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][205]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][206]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][206]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][206] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][206]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][207]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][207]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][207] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][207]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][208]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][208]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][208] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][208]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][209]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][209]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][209] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][209]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][20]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][20]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][20] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][20]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][210]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][210]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][210] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][210]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][211]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][211]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][211] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][211]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][212]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][212]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][212] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][212]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][213]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][213]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][213] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][213]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][214]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][214]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][214] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][214]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][215]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][215]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][215] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][215]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][216]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][216]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][216] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][216]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][217]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][217]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][217] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][217]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][218]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][218]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][218] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][218]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][219]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][219]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][219] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][219]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][21]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][21]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][21] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][21]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][220]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][220]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][220] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][220]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][221]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][221]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][221] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][221]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][222]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][222]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][222] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][222]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][223]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][223]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][223] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][223]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][224]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][224]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][224] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][224]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][225]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][225]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][225] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][225]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][226]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][226]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][226] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][226]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][227]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][227]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][227] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][227]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][228]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][228]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][228] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][228]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][229]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][229]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][229] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][229]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][22]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][22]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][22] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][22]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][230]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][230]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][230] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][230]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][231]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][231]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][231] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][231]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][232]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][232]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][232] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][232]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][233]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][233]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][233] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][233]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][234]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][234]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][234] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][234]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][235]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][235]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][235] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][235]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][236]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][236]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][236] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][236]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][237]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][237]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][237] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][237]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][238]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][238]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][238] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][238]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][239]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][239]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][239] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][239]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][23]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][23]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][23] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][23]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][240]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][240]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][240] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][240]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][241]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][241]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][241] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][241]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][242]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][242]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][242] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][242]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][243]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][243]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][243] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][243]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][244]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][244]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][244] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][244]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][245]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][245]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][245] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][245]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][246]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][246]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][246] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][246]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][247]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][247]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][247] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][247]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][248]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][248]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][248] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][248]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][249]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][249]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][249] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][249]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][24]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][24]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][24] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][24]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][250]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][250]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][250] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][250]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][251]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][251]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][251] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][251]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][252]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][252]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][252] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][252]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][253]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][253]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][253] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][253]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][254]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][254]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][254] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][254]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][255]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][255]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][255] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][255]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][256]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][256]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][256] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][256]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][257]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][257]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][257] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][257]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][258]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][258]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][258] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][258]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][259]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][259]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][259] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][259]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][25]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][25]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][25] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][25]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][260]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][260]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][260] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][260]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][261]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][261]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][261] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][261]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][262]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][262]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][262] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][262]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][263]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][263]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][263] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][263]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][264]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][264]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][264] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][264]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][265]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][265]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][265] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][265]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][266]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][266]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][266] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][266]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][267]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][267]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][267] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][267]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][268]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][268]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][268] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][268]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][269]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][269]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][269] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][269]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][26]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][26]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][26] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][26]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][270]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][270]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][270] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][270]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][271]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][271]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][271] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][271]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][272]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][272]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][272] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][272]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][273]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][273]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][273] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][273]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][274]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][274]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][274] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][274]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][275]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][275]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][275] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][275]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][276]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][276]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][276] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][276]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][277]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][277]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][277] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][277]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][278]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][278]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][278] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][278]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][279]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][279]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][279] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][279]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][27]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][27]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][27] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][27]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][280]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][280]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][280] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][280]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][281]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][281]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][281] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][281]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][282]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][282]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][282] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][282]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][283]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][283]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][283] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][283]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][284]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][284]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][284] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][284]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][285]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][285]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][285] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][285]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][286]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][286]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][286] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][286]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][287]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][287]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][287] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][287]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][288]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][288]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][288] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][288]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][289]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][289]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][289] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][289]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][28]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][28]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][28] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][28]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][290]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][290]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][290] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][290]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][291]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][291]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][291] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][291]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][292]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][292]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][292] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][292]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][293]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][293]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][293] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][293]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][294]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][294]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][294] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][294]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][295]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][295]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][295] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][295]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][296]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][296]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][296] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][296]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][297]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][297]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][297] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][297]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][298]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][298]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][298] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][298]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][299]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][299]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][299] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][299]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][29]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][29]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][29] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][29]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][2]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][2]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][2] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][2]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][300]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][300]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][300] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][300]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][301]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][301]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][301] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][301]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][302]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][302]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][302] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][302]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][303]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][303]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][303] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][303]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][304]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][304]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][304] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][304]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][305]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][305]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][305] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][305]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][306]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][306]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][306] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][306]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][307]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][307]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][307] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][307]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][308]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][308]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][308] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][308]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][309]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][309]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][309] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][309]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][30]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][30]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][30] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][30]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][310]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][310]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][310] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][310]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][311]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][311]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][311] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][311]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][312]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][312]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][312] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][312]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][313]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][313]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][313] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][313]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][314]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][314]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][314] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][314]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][315]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][315]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][315] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][315]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][316]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][316]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][316] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][316]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][317]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][317]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][317] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][317]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][318]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][318]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][318] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][318]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][319]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][319]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][319] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][319]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][31]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][31]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][31] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][31]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][320]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][320]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][320] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][320]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][321]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][321]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][321] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][321]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][322]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][322]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][322] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][322]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][323]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][323]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][323] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][323]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][324]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][324]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][324] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][324]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][325]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][325]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][325] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][325]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][326]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][326]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][326] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][326]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][327]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][327]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][327] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][327]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][328]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][328]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][328] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][328]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][329]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][329]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][329] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][329]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][32]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][32]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][32] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][32]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][330]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][330]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][330] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][330]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][331]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][331]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][331] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][331]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][332]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][332]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][332] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][332]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][333]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][333]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][333] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][333]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][334]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][334]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][334] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][334]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][335]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][335]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][335] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][335]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][336]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][336]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][336] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][336]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][337]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][337]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][337] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][337]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][338]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][338]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][338] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][338]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][339]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][339]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][339] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][339]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][33]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][33]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][33] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][33]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][340]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][340]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][340] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][340]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][341]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][341]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][341] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][341]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][342]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][342]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][342] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][342]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][343]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][343]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][343] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][343]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][344]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][344]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][344] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][344]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][345]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][345]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][345] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][345]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][346]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][346]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][346] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][346]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][347]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][347]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][347] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][347]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][348]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][348]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][348] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][348]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][349]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][349]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][349] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][349]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][34]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][34]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][34] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][34]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][350]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][350]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][350] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][350]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][351]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][351]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][351] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][351]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][352]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][352]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][352] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][352]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][353]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][353]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][353] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][353]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][354]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][354]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][354] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][354]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][355]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][355]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][355] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][355]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][356]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][356]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][356] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][356]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][357]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][357]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][357] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][357]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][358]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][358]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][358] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][358]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][359]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][359]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][359] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][359]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][35]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][35]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][35] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][35]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][360]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][360]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][360] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][360]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][361]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][361]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][361] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][361]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][362]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][362]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][362] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][362]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][363]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][363]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][363] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][363]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][364]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][364]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][364] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][364]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][365]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][365]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][365] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][365]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][366]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][366]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][366] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][366]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][367]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][367]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][367] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][367]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][368]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][368]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][368] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][368]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][369]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][369]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][369] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][369]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][36]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][36]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][36] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][36]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][370]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][370]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][370] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][370]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][371]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][371]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][371] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][371]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][372]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][372]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][372] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][372]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][373]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][373]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][373] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][373]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][374]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][374]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][374] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][374]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][375]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][375]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][375] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][375]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][376]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][376]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][376] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][376]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][377]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][377]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][377] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][377]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][378]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][378]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][378] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][378]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][379]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][379]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][379] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][379]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][37]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][37]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][37] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][37]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][380]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][380]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][380] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][380]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][381]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][381]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][381] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][381]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][382]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][382]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][382] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][382]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][383]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][383]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][383] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][383]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][384]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][384]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][384] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][384]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][385]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][385]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][385] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][385]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][386]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][386]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][386] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][386]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][387]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][387]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][387] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][387]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][388]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][388]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][388] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][388]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][389]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][389]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][389] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][389]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][38]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][38]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][38] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][38]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][390]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][390]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][390] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][390]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][391]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][391]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][391] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][391]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][392]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][392]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][392] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][392]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][393]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][393]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][393] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][393]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][394]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][394]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][394] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][394]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][395]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][395]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][395] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][395]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][396]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][396]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][396] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][396]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][397]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][397]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][397] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][397]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][398]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][398]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][398] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][398]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][399]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][399]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][399] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][399]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][39]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][39]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][39] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][39]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][3]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][3]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][3] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][3]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][400]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][400]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][400] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][400]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][401]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][401]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][401] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][401]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][402]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][402]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][402] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][402]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][403]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][403]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][403] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][403]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][404]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][404]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][404] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][404]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][405]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][405]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][405] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][405]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][406]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][406]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][406] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][406]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][407]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][407]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][407] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][407]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][408]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][408]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][408] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][408]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][409]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][409]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][409] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][409]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][40]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][40]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][40] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][40]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][410]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][410]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][410] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][410]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][411]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][411]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][411] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][411]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][412]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][412]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][412] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][412]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][413]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][413]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][413] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][413]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][414]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][414]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][414] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][414]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][415]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][415]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][415] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][415]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][416]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][416]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][416] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][416]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][417]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][417]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][417] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][417]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][418]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][418]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][418] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][418]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][419]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][419]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][419] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][419]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][41]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][41]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][41] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][41]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][420]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][420]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][420] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][420]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][421]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][421]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][421] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][421]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][422]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][422]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][422] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][422]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][423]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][423]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][423] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][423]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][424]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][424]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][424] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][424]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][425]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][425]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][425] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][425]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][426]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][426]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][426] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][426]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][427]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][427]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][427] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][427]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][428]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][428]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][428] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][428]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][429]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][429]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][429] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][429]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][42]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][42]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][42] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][42]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][430]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][430]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][430] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][430]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][431]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][431]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][431] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][431]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][432]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][432]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][432] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][432]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][433]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][433]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][433] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][433]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][434]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][434]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][434] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][434]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][435]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][435]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][435] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][435]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][436]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][436]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][436] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][436]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][437]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][437]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][437] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][437]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][438]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][438]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][438] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][438]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][439]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][439]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][439] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][439]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][43]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][43]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][43] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][43]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][440]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][440]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][440] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][440]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][441]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][441]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][441] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][441]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][442]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][442]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][442] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][442]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][443]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][443]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][443] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][443]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][444]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][444]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][444] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][444]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][445]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][445]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][445] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][445]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][446]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][446]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][446] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][446]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][447]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][447]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][447] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][447]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][448]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][448]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][448] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][448]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][449]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][449]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][449] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][449]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][44]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][44]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][44] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][44]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][450]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][450]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][450] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][450]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][451]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][451]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][451] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][451]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][452]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][452]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][452] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][452]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][453]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][453]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][453] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][453]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][454]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][454]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][454] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][454]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][455]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][455]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][455] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][455]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][456]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][456]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][456] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][456]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][457]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][457]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][457] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][457]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][458]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][458]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][458] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][458]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][459]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][459]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][459] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][459]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][45]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][45]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][45] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][45]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][460]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][460]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][460] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][460]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][461]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][461]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][461] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][461]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][462]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][462]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][462] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][462]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][463]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][463]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][463] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][463]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][464]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][464]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][464] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][464]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][465]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][465]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][465] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][465]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][466]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][466]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][466] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][466]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][467]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][467]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][467] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][467]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][468]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][468]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][468] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][468]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][469]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][469]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][469] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][469]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][46]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][46]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][46] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][46]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][470]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][470]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][470] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][470]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][471]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][471]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][471] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][471]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][472]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][472]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][472] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][472]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][473]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][473]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][473] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][473]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][474]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][474]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][474] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][474]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][475]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][475]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][475] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][475]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][476]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][476]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][476] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][476]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][477]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][477]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][477] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][477]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][478]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][478]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][478] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][478]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][479]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][479]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][479] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][479]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][47]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][47]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][47] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][47]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][480]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][480]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][480] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][480]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][481]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][481]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][481] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][481]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][482]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][482]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][482] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][482]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][483]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][483]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][483] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][483]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][484]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][484]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][484] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][484]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][485]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][485]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][485] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][485]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][486]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][486]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][486] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][486]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][487]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][487]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][487] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][487]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][488]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][488]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][488] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][488]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][489]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][489]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][489] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][489]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][48]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][48]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][48] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][48]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][490]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][490]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][490] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][490]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][491]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][491]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][491] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][491]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][492]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][492]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][492] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][492]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][493]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][493]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][493] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][493]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][494]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][494]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][494] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][494]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][495]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][495]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][495] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][495]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][496]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][496]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][496] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][496]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][497]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][497]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][497] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][497]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][498]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][498]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][498] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][498]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][499]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][499]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][499] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][499]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][49]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][49]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][49] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][49]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][4]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][4]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][4] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][4]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][500]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][500]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][500] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][500]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][501]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][501]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][501] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][501]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][502]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][502]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][502] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][502]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][503]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][503]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][503] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][503]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][504]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][504]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][504] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][504]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][505]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][505]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][505] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][505]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][506]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][506]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][506] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][506]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][507]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][507]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][507] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][507]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][508]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][508]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][508] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][508]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][509]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][509]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][509] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][509]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][50]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][50]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][50] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][50]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][510]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][510]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][510] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][510]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][511]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][511]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][511] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][511]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][512]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][512]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][512] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][512]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][513]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][513]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][513] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][513]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][514]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][514]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][514] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][514]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][515]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][515]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][515] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][515]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][516]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][516]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][516] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][516]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][517]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][517]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][517] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][517]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][518]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][518]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][518] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][518]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][519]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][519]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][519] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][519]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][51]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][51]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][51] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][51]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][520]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][520]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][520] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][520]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][521]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][521]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][521] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][521]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][522]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][522]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][522] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][522]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][523]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][523]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][523] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][523]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][524]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][524]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][524] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][524]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][525]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][525]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][525] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][525]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][526]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][526]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][526] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][526]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][527]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][527]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][527] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][527]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][528]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][528]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][528] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][528]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][529]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][529]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][529] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][529]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][52]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][52]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][52] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][52]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][530]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][530]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][530] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][530]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][531]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][531]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][531] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][531]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][532]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][532]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][532] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][532]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][533]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][533]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][533] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][533]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][534]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][534]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][534] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][534]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][535]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][535]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][535] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][535]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][536]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][536]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][536] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][536]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][537]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][537]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][537] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][537]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][538]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][538]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][538] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][538]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][539]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][539]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][539] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][539]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][53]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][53]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][53] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][53]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][540]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][540]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][540] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][540]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][541]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][541]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][541] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][541]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][542]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][542]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][542] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][542]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][543]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][543]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][543] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][543]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][544]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][544]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][544] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][544]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][545]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][545]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][545] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][545]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][546]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][546]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][546] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][546]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][547]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][547]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][547] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][547]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][548]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][548]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][548] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][548]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][549]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][549]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][549] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][549]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][54]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][54]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][54] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][54]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][550]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][550]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][550] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][550]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][551]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][551]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][551] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][551]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][552]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][552]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][552] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][552]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][553]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][553]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][553] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][553]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][554]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][554]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][554] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][554]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][555]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][555]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][555] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][555]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][556]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][556]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][556] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][556]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][557]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][557]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][557] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][557]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][558]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][558]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][558] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][558]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][559]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][559]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][559] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][559]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][55]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][55]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][55] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][55]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][560]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][560]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][560] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][560]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][561]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][561]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][561] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][561]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][562]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][562]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][562] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][562]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][563]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][563]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][563] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][563]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][564]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][564]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][564] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][564]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][565]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][565]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][565] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][565]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][566]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][566]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][566] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][566]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][567]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][567]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][567] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][567]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][568]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][568]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][568] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][568]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][569]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][569]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][569] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][569]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][56]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][56]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][56] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][56]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][570]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][570]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][570] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][570]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][571]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][571]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][571] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][571]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][572]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][572]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][572] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][572]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][573]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][573]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][573] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][573]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][574]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][574]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][574] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][574]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][575]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][575]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][575] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][575]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][576]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][576]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][576] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][576]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][577]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][577]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][577] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][577]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][578]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][578]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][578] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][578]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][579]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][579]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][579] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][579]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][57]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][57]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][57] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][57]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][580]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][580]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][580] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][580]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][581]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][581]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][581] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][581]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][582]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][582]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][582] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][582]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][583]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][583]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][583] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][583]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][584]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][584]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][584] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][584]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][585]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][585]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][585] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][585]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][586]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][586]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][586] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][586]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][587]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][587]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][587] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][587]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][588]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][588]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][588] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][588]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][589]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][589]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][589] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][589]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][58]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][58]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][58] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][58]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][590]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][590]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][590] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][590]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][591]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][591]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][591] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][591]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][592]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][592]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][592] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][592]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][593]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][593]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][593] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][593]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][594]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][594]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][594] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][594]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][595]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][595]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][595] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][595]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][596]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][596]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][596] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][596]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][597]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][597]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][597] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][597]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][598]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][598]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][598] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][598]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][599]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][599]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][599] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][599]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][59]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][59]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][59] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][59]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][5]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][5]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][5] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][5]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][600]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][600]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][600] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][600]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][601]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][601]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][601] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][601]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][602]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][602]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][602] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][602]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][603]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][603]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][603] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][603]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][604]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][604]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][604] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][604]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][605]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][605]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][605] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][605]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][606]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][606]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][606] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][606]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][607]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][607]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][607] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][607]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][608]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][608]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][608] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][608]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][609]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][609]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][609] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][609]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][60]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][60]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][60] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][60]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][610]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][610]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][610] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][610]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][611]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][611]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][611] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][611]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][612]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][612]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][612] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][612]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][613]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][613]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][613] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][613]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][614]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][614]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][614] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][614]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][615]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][615]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][615] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][615]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][616]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][616]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][616] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][616]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][617]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][617]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][617] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][617]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][618]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][618]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][618] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][618]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][619]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][619]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][619] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][619]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][61]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][61]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][61] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][61]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][620]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][620]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][620] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][620]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][621]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][621]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][621] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][621]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][622]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][622]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][622] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][622]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][623]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][623]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][623] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][623]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][624]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][624]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][624] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][624]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][625]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][625]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][625] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][625]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][626]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][626]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][626] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][626]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][627]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][627]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][627] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][627]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][628]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][628]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][628] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][628]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][629]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][629]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][629] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][629]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][62]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][62]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][62] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][62]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][630]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][630]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][630] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][630]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][631]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][631]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][631] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][631]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][632]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][632]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][632] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][632]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][633]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][633]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][633] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][633]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][634]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][634]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][634] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][634]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][635]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][635]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][635] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][635]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][636]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][636]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][636] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][636]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][637]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][637]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][637] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][637]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][638]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][638]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][638] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][638]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][639]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][639]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][639] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][639]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][63]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][63]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][63] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][63]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][640]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][640]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][640] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][640]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][641]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][641]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][641] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][641]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][642]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][642]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][642] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][642]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][643]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][643]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][643] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][643]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][644]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][644]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][644] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][644]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][645]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][645]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][645] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][645]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][646]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][646]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][646] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][646]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][647]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][647]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][647] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][647]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][648]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][648]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][648] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][648]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][649]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][649]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][649] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][649]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][64]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][64]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][64] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][64]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][650]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][650]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][650] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][650]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][651]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][651]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][651] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][651]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][652]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][652]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][652] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][652]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][653]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][653]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][653] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][653]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][654]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][654]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][654] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][654]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][655]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][655]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][655] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][655]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][656]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][656]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][656] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][656]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][657]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][657]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][657] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][657]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][658]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][658]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][658] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][658]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][659]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][659]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][659] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][659]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][65]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][65]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][65] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][65]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][660]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][660]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][660] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][660]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][661]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][661]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][661] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][661]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][662]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][662]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][662] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][662]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][663]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][663]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][663] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][663]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][664]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][664]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][664] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][664]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][665]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][665]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][665] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][665]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][666]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][666]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][666] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][666]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][667]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][667]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][667] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][667]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][668]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][668]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][668] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][668]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][669]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][669]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][669] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][669]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][66]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][66]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][66] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][66]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][670]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][670]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][670] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][670]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][671]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][671]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][671] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][671]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][672]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][672]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][672] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][672]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][673]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][673]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][673] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][673]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][674]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][674]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][674] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][674]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][675]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][675]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][675] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][675]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][676]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][676]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][676] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][676]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][677]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][677]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][677] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][677]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][678]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][678]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][678] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][678]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][679]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][679]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][679] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][679]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][67]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][67]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][67] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][67]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][680]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][680]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][680] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][680]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][681]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][681]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][681] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][681]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][682]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][682]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][682] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][682]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][683]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][683]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][683] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][683]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][684]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][684]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][684] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][684]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][685]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][685]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][685] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][685]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][686]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][686]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][686] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][686]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][687]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][687]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][687] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][687]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][688]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][688]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][688] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][688]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][689]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][689]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][689] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][689]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][68]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][68]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][68] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][68]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][690]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][690]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][690] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][690]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][691]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][691]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][691] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][691]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][692]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][692]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][692] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][692]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][693]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][693]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][693] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][693]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][694]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][694]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][694] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][694]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][695]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][695]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][695] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][695]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][696]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][696]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][696] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][696]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][697]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][697]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][697] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][697]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][698]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][698]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][698] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][698]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][699]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][699]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][699] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][699]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][69]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][69]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][69] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][69]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][6]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][6]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][6] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][6]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][700]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][700]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][700] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][700]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][701]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][701]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][701] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][701]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][702]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][702]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][702] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][702]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][703]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][703]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][703] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][703]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][704]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][704]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][704] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][704]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][705]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][705]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][705] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][705]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][706]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][706]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][706] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][706]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][707]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][707]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][707] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][707]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][708]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][708]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][708] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][708]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][709]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][709]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][709] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][709]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][70]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][70]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][70] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][70]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][710]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][710]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][710] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][710]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][711]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][711]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][711] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][711]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][712]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][712]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][712] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][712]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][713]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][713]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][713] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][713]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][714]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][714]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][714] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][714]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][715]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][715]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][715] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][715]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][716]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][716]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][716] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][716]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][717]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][717]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][717] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][717]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][718]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][718]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][718] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][718]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][719]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][719]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][719] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][719]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][71]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][71]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][71] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][71]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][720]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][720]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][720] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][720]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][721]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][721]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][721] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][721]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][722]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][722]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][722] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][722]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][723]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][723]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][723] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][723]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][724]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][724]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][724] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][724]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][725]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][725]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][725] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][725]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][726]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][726]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][726] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][726]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][727]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][727]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][727] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][727]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][728]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][728]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][728] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][728]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][729]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][729]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][729] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][729]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][72]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][72]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][72] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][72]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][730]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][730]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][730] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][730]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][731]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][731]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][731] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][731]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][732]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][732]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][732] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][732]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][733]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][733]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][733] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][733]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][734]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][734]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][734] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][734]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][735]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][735]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][735] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][735]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][736]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][736]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][736] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][736]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][737]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][737]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][737] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][737]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][738]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][738]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][738] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][738]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][739]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][739]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][739] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][739]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][73]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][73]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][73] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][73]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][740]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][740]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][740] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][740]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][741]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][741]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][741] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][741]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][742]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][742]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][742] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][742]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][743]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][743]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][743] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][743]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][744]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][744]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][744] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][744]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][745]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][745]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][745] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][745]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][746]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][746]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][746] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][746]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][747]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][747]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][747] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][747]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][748]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][748]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][748] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][748]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][749]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][749]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][749] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][749]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][74]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][74]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][74] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][74]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][750]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][750]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][750] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][750]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][751]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][751]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][751] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][751]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][752]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][752]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][752] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][752]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][753]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][753]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][753] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][753]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][754]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][754]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][754] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][754]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][755]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][755]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][755] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][755]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][756]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][756]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][756] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][756]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][757]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][757]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][757] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][757]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][758]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][758]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][758] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][758]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][759]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][759]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][759] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][759]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][75]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][75]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][75] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][75]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][760]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][760]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][760] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][760]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][761]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][761]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][761] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][761]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][762]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][762]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][762] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][762]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][763]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][763]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][763] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][763]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][764]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][764]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][764] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][764]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][765]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][765]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][765] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][765]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][766]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][766]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][766] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][766]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][767]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][767]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][767] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][767]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][768]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][768]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][768] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][768]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][769]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][769]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][769] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][769]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][76]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][76]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][76] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][76]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][770]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][770]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][770] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][770]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][771]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][771]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][771] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][771]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][772]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][772]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][772] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][772]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][773]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][773]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][773] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][773]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][774]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][774]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][774] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][774]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][775]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][775]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][775] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][775]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][776]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][776]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][776] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][776]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][777]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][777]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][777] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][777]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][778]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][778]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][778] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][778]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][779]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][779]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][779] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][779]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][77]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][77]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][77] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][77]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][780]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][780]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][780] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][780]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][781]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][781]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][781] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][781]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][782]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][782]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][782] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][782]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][783]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][783]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][783] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][783]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][784]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][784]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][784] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][784]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][785]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][785]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][785] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][785]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][786]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][786]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][786] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][786]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][787]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][787]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][787] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][787]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][788]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][788]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][788] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][788]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][789]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][789]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][789] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][789]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][78]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][78]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][78] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][78]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][790]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][790]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][790] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][790]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][791]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][791]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][791] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][791]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][792]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][792]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][792] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][792]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][793]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][793]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][793] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][793]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][794]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][794]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][794] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][794]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][795]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][795]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][795] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][795]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][796]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][796]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][796] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][796]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][797]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][797]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][797] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][797]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][798]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][798]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][798] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][798]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][799]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][799]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][799] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][799]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][79]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][79]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][79] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][79]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][7]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][7]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][7] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][7]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][800]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][800]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][800] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][800]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][801]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][801]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][801] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][801]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][802]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][802]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][802] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][802]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][803]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][803]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][803] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][803]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][804]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][804]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][804] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][804]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][805]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][805]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][805] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][805]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][806]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][806]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][806] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][806]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][807]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][807]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][807] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][807]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][808]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][808]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][808] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][808]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][809]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][809]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][809] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][809]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][80]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][80]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][80] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][80]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][810]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][810]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][810] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][810]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][811]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][811]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][811] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][811]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][812]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][812]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][812] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][812]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][813]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][813]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][813] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][813]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][814]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][814]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][814] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][814]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][815]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][815]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][815] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][815]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][816]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][816]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][816] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][816]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][817]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][817]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][817] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][817]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][818]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][818]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][818] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][818]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][819]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][819]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][819] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][819]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][81]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][81]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][81] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][81]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][820]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][820]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][820] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][820]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][821]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][821]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][821] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][821]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][822]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][822]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][822] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][822]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][823]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][823]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][823] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][823]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][824]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][824]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][824] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][824]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][825]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][825]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][825] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][825]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][826]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][826]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][826] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][826]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][827]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][827]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][827] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][827]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][828]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][828]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][828] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][828]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][829]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][829]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][829] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][829]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][82]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][82]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][82] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][82]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][830]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][830]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][830] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][830]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][831]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][831]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][831] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][831]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][832]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][832]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][832] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][832]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][833]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][833]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][833] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][833]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][834]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][834]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][834] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][834]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][835]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][835]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][835] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][835]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][836]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][836]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][836] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][836]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][837]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][837]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][837] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][837]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][838]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][838]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][838] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][838]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][839]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][839]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][839] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][839]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][83]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][83]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][83] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][83]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][840]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][840]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][840] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][840]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][841]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][841]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][841] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][841]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][842]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][842]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][842] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][842]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][843]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][843]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][843] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][843]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][844]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][844]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][844] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][844]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][845]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][845]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][845] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][845]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][846]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][846]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][846] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][846]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][847]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][847]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][847] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][847]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][848]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][848]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][848] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][848]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][849]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][849]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][849] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][849]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][84]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][84]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][84] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][84]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][850]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][850]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][850] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][850]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][851]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][851]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][851] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][851]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][852]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][852]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][852] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][852]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][853]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][853]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][853] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][853]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][854]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][854]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][854] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][854]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][855]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][855]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][855] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][855]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][856]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][856]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][856] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][856]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][857]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][857]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][857] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][857]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][858]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][858]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][858] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][858]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][859]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][859]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][859] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][859]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][85]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][85]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][85] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][85]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][860]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][860]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][860] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][860]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][861]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][861]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][861] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][861]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][862]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][862]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][862] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][862]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][863]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][863]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][863] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][863]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][864]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][864]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][864] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][864]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][865]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][865]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][865] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][865]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][866]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][866]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][866] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][866]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][867]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][867]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][867] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][867]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][868]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][868]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][868] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][868]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][869]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][869]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][869] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][869]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][86]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][86]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][86] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][86]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][870]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][870]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][870] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][870]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][871]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][871]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][871] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][871]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][872]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][872]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][872] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][872]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][873]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][873]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][873] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][873]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][874]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][874]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][874] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][874]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][875]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][875]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][875] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][875]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][876]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][876]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][876] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][876]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][877]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][877]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][877] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][877]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][878]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][878]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][878] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][878]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][879]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][879]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][879] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][879]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][87]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][87]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][87] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][87]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][880]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][880]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][880] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][880]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][881]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][881]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][881] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][881]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][882]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][882]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][882] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][882]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][883]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][883]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][883] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][883]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][884]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][884]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][884] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][884]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][885]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][885]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][885] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][885]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][886]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][886]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][886] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][886]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][887]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][887]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][887] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][887]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][888]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][888]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][888] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][888]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][889]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][889]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][889] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][889]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][88]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][88]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][88] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][88]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][890]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][890]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][890] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][890]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][891]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][891]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][891] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][891]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][892]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][892]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][892] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][892]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][893]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][893]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][893] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][893]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][894]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][894]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][894] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][894]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][895]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][895]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][895] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][895]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][896]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][896]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][896] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][896]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][897]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][897]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][897] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][897]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][898]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][898]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][898] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][898]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][899]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][899]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][899] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][899]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][89]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][89]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][89] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][89]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][8]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][8]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][8] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][8]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][900]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][900]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][900] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][900]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][901]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][901]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][901] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][901]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][902]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][902]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][902] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][902]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][903]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][903]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][903] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][903]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][904]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][904]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][904] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][904]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][905]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][905]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][905] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][905]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][906]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][906]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][906] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][906]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][907]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][907]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][907] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][907]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][908]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][908]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][908] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][908]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][909]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][909]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][909] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][909]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][90]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][90]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][90] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][90]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][910]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][910]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][910] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][910]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][911]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][911]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][911] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][911]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][912]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][912]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][912] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][912]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][913]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][913]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][913] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][913]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][914]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][914]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][914] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][914]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][915]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][915]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][915] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][915]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][916]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][916]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][916] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][916]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][917]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][917]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][917] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][917]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][918]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][918]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][918] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][918]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][919]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][919]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][919] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][919]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][91]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][91]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][91] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][91]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][920]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][920]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][920] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][920]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][921]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][921]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][921] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][921]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][922]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][922]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][922] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][922]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][923]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][923]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][923] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][923]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][924]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][924]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][924] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][924]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][925]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][925]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][925] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][925]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][926]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][926]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][926] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][926]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][927]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][927]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][927] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][927]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][928]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][928]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][928] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][928]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][929]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][929]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][929] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][929]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][92]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][92]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][92] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][92]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][930]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][930]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][930] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][930]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][931]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][931]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][931] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][931]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][932]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][932]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][932] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][932]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][933]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][933]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][933] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][933]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][934]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][934]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][934] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][934]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][935]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][935]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][935] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][935]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][936]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][936]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][936] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][936]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][937]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][937]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][937] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][937]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][938]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][938]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][938] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][938]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][939]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][939]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][939] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][939]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][93]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][93]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][93] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][93]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][940]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][940]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][940] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][940]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][941]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][941]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][941] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][941]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][942]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][942]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][942] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][942]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][943]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][943]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][943] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][943]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][944]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][944]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][944] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][944]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][945]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][945]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][945] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][945]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][946]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][946]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][946] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][946]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][947]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][947]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][947] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][947]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][948]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][948]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][948] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][948]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][949]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][949]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][949] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][949]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][94]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][94]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][94] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][94]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][950]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][950]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][950] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][950]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][951]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][951]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][951] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][951]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][952]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][952]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][952] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][952]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][953]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][953]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][953] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][953]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][954]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][954]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][954] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][954]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][955]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][955]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][955] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][955]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][956]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][956]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][956] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][956]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][957]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][957]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][957] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][957]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][958]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][958]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][958] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][958]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][959]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][959]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][959] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][959]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][95]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][95]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][95] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][95]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][960]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][960]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][960] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][960]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][961]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][961]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][961] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][961]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][962]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][962]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][962] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][962]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][963]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][963]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][963] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][963]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][964]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][964]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][964] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][964]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][965]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][965]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][965] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][965]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][966]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][966]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][966] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][966]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][967]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][967]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][967] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][967]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][968]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][968]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][968] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][968]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][969]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][969]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][969] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][969]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][96]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][96]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][96] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][96]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][970]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][970]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][970] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][970]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][971]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][971]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][971] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][971]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][972]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][972]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][972] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][972]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][973]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][973]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][973] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][973]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][974]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][974]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][974] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][974]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][975]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][975]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][975] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][975]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][976]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][976]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][976] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][976]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][977]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][977]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][977] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][977]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][978]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][978]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][978] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][978]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][979]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][979]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][979] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][979]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][97]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][97]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][97] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][97]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][980]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][980]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][980] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][980]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][981]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][981]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][981] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][981]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][982]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][982]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][982] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][982]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][983]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][983]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][983] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][983]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][984]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][984]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][984] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][984]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][985]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][985]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][985] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][985]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][986]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][986]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][986] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][986]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][987]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][987]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][987] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][987]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][988]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][988]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][988] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][988]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][989]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][989]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][989] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][989]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][98]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][98]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][98] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][98]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][990]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][990]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][990] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][990]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][991]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][991]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][991] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][991]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][992]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][992]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][992] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][992]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][993]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][993]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][993] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][993]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][994]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][994]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][994] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][994]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][995]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][995]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][995] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][995]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][996]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][996]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][996] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][996]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][997]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][997]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][997] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][997]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][998]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][998]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][998] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][998]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][999]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][999]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][999] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][999]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][99]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][99]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][99] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][99]_srl3_n_0 ));
  (* srl_bus_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4] " *) 
  (* srl_name = "\\i_shiftreg_point/DELAY_BLOCK[3].shift_array_reg[4][9]_srl3 " *) 
  SRL16E #(
    .INIT(16'h0000)) 
    \DELAY_BLOCK[3].shift_array_reg[4][9]_srl3 
       (.A0(\<const0> ),
        .A1(\<const1> ),
        .A2(\<const0> ),
        .A3(\<const0> ),
        .CE(\<const1> ),
        .CLK(clk),
        .D(\shift_array_reg_n_0_[1][9] ),
        .Q(\DELAY_BLOCK[3].shift_array_reg[4][9]_srl3_n_0 ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][0]_srl3_n_0 ),
        .Q(acc_point_o[0]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1000] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1000]_srl3_n_0 ),
        .Q(acc_point_o[1000]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1001] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1001]_srl3_n_0 ),
        .Q(acc_point_o[1001]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1002] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1002]_srl3_n_0 ),
        .Q(acc_point_o[1002]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1003] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1003]_srl3_n_0 ),
        .Q(acc_point_o[1003]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1004] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1004]_srl3_n_0 ),
        .Q(acc_point_o[1004]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1005] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1005]_srl3_n_0 ),
        .Q(acc_point_o[1005]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1006] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1006]_srl3_n_0 ),
        .Q(acc_point_o[1006]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1007] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1007]_srl3_n_0 ),
        .Q(acc_point_o[1007]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1008] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1008]_srl3_n_0 ),
        .Q(acc_point_o[1008]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1009] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1009]_srl3_n_0 ),
        .Q(acc_point_o[1009]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][100] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][100]_srl3_n_0 ),
        .Q(acc_point_o[100]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1010] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1010]_srl3_n_0 ),
        .Q(acc_point_o[1010]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1011] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1011]_srl3_n_0 ),
        .Q(acc_point_o[1011]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1012] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1012]_srl3_n_0 ),
        .Q(acc_point_o[1012]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1013] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1013]_srl3_n_0 ),
        .Q(acc_point_o[1013]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1014] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1014]_srl3_n_0 ),
        .Q(acc_point_o[1014]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1015] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1015]_srl3_n_0 ),
        .Q(acc_point_o[1015]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1016] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1016]_srl3_n_0 ),
        .Q(acc_point_o[1016]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1017] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1017]_srl3_n_0 ),
        .Q(acc_point_o[1017]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1018] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1018]_srl3_n_0 ),
        .Q(acc_point_o[1018]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1019] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1019]_srl3_n_0 ),
        .Q(acc_point_o[1019]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][101] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][101]_srl3_n_0 ),
        .Q(acc_point_o[101]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1020] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1020]_srl3_n_0 ),
        .Q(acc_point_o[1020]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1021] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1021]_srl3_n_0 ),
        .Q(acc_point_o[1021]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1022] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1022]_srl3_n_0 ),
        .Q(acc_point_o[1022]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1023] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1023]_srl3_n_0 ),
        .Q(acc_point_o[1023]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1024] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1024]_srl3_n_0 ),
        .Q(acc_point_o[1024]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1025] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1025]_srl3_n_0 ),
        .Q(acc_point_o[1025]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1026] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1026]_srl3_n_0 ),
        .Q(acc_point_o[1026]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1027] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1027]_srl3_n_0 ),
        .Q(acc_point_o[1027]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1028] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1028]_srl3_n_0 ),
        .Q(acc_point_o[1028]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1029] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1029]_srl3_n_0 ),
        .Q(acc_point_o[1029]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][102] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][102]_srl3_n_0 ),
        .Q(acc_point_o[102]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1030] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1030]_srl3_n_0 ),
        .Q(acc_point_o[1030]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1031] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1031]_srl3_n_0 ),
        .Q(acc_point_o[1031]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1032] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1032]_srl3_n_0 ),
        .Q(acc_point_o[1032]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1033] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1033]_srl3_n_0 ),
        .Q(acc_point_o[1033]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1034] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1034]_srl3_n_0 ),
        .Q(acc_point_o[1034]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1035] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1035]_srl3_n_0 ),
        .Q(acc_point_o[1035]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1036] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1036]_srl3_n_0 ),
        .Q(acc_point_o[1036]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1037] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1037]_srl3_n_0 ),
        .Q(acc_point_o[1037]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1038] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1038]_srl3_n_0 ),
        .Q(acc_point_o[1038]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1039] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1039]_srl3_n_0 ),
        .Q(acc_point_o[1039]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][103] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][103]_srl3_n_0 ),
        .Q(acc_point_o[103]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1040] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1040]_srl3_n_0 ),
        .Q(acc_point_o[1040]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1041] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1041]_srl3_n_0 ),
        .Q(acc_point_o[1041]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1042] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1042]_srl3_n_0 ),
        .Q(acc_point_o[1042]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1043] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1043]_srl3_n_0 ),
        .Q(acc_point_o[1043]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1044] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1044]_srl3_n_0 ),
        .Q(acc_point_o[1044]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1045] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1045]_srl3_n_0 ),
        .Q(acc_point_o[1045]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1046] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1046]_srl3_n_0 ),
        .Q(acc_point_o[1046]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1047] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1047]_srl3_n_0 ),
        .Q(acc_point_o[1047]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1048] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1048]_srl3_n_0 ),
        .Q(acc_point_o[1048]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1049] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1049]_srl3_n_0 ),
        .Q(acc_point_o[1049]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][104] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][104]_srl3_n_0 ),
        .Q(acc_point_o[104]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1050] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1050]_srl3_n_0 ),
        .Q(acc_point_o[1050]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1051] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1051]_srl3_n_0 ),
        .Q(acc_point_o[1051]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1052] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1052]_srl3_n_0 ),
        .Q(acc_point_o[1052]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1053] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1053]_srl3_n_0 ),
        .Q(acc_point_o[1053]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1054] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1054]_srl3_n_0 ),
        .Q(acc_point_o[1054]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1055] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1055]_srl3_n_0 ),
        .Q(acc_point_o[1055]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1056] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1056]_srl3_n_0 ),
        .Q(acc_point_o[1056]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1057] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1057]_srl3_n_0 ),
        .Q(acc_point_o[1057]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1058] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1058]_srl3_n_0 ),
        .Q(acc_point_o[1058]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1059] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1059]_srl3_n_0 ),
        .Q(acc_point_o[1059]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][105] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][105]_srl3_n_0 ),
        .Q(acc_point_o[105]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1060] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1060]_srl3_n_0 ),
        .Q(acc_point_o[1060]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1061] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1061]_srl3_n_0 ),
        .Q(acc_point_o[1061]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1062] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1062]_srl3_n_0 ),
        .Q(acc_point_o[1062]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1063] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1063]_srl3_n_0 ),
        .Q(acc_point_o[1063]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1064] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1064]_srl3_n_0 ),
        .Q(acc_point_o[1064]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1065] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1065]_srl3_n_0 ),
        .Q(acc_point_o[1065]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1066] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1066]_srl3_n_0 ),
        .Q(acc_point_o[1066]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1067] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1067]_srl3_n_0 ),
        .Q(acc_point_o[1067]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1068] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1068]_srl3_n_0 ),
        .Q(acc_point_o[1068]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1069] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1069]_srl3_n_0 ),
        .Q(acc_point_o[1069]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][106] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][106]_srl3_n_0 ),
        .Q(acc_point_o[106]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1070] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1070]_srl3_n_0 ),
        .Q(acc_point_o[1070]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1071] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1071]_srl3_n_0 ),
        .Q(acc_point_o[1071]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1072] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1072]_srl3_n_0 ),
        .Q(acc_point_o[1072]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1073] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1073]_srl3_n_0 ),
        .Q(acc_point_o[1073]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1074] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1074]_srl3_n_0 ),
        .Q(acc_point_o[1074]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1075] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1075]_srl3_n_0 ),
        .Q(acc_point_o[1075]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1076] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1076]_srl3_n_0 ),
        .Q(acc_point_o[1076]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1077] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1077]_srl3_n_0 ),
        .Q(acc_point_o[1077]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1078] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1078]_srl3_n_0 ),
        .Q(acc_point_o[1078]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1079] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1079]_srl3_n_0 ),
        .Q(acc_point_o[1079]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][107] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][107]_srl3_n_0 ),
        .Q(acc_point_o[107]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1080] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1080]_srl3_n_0 ),
        .Q(acc_point_o[1080]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1081] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1081]_srl3_n_0 ),
        .Q(acc_point_o[1081]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1082] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1082]_srl3_n_0 ),
        .Q(acc_point_o[1082]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1083] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1083]_srl3_n_0 ),
        .Q(acc_point_o[1083]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1084] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1084]_srl3_n_0 ),
        .Q(acc_point_o[1084]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1085] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1085]_srl3_n_0 ),
        .Q(acc_point_o[1085]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1086] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1086]_srl3_n_0 ),
        .Q(acc_point_o[1086]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1087] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1087]_srl3_n_0 ),
        .Q(acc_point_o[1087]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1088] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1088]_srl3_n_0 ),
        .Q(acc_point_o[1088]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1089] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1089]_srl3_n_0 ),
        .Q(acc_point_o[1089]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][108] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][108]_srl3_n_0 ),
        .Q(acc_point_o[108]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1090] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1090]_srl3_n_0 ),
        .Q(acc_point_o[1090]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1091] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1091]_srl3_n_0 ),
        .Q(acc_point_o[1091]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1092] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1092]_srl3_n_0 ),
        .Q(acc_point_o[1092]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1093] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1093]_srl3_n_0 ),
        .Q(acc_point_o[1093]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1094] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1094]_srl3_n_0 ),
        .Q(acc_point_o[1094]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1095] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1095]_srl3_n_0 ),
        .Q(acc_point_o[1095]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1096] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1096]_srl3_n_0 ),
        .Q(acc_point_o[1096]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1097] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1097]_srl3_n_0 ),
        .Q(acc_point_o[1097]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1098] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1098]_srl3_n_0 ),
        .Q(acc_point_o[1098]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1099] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1099]_srl3_n_0 ),
        .Q(acc_point_o[1099]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][109] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][109]_srl3_n_0 ),
        .Q(acc_point_o[109]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][10]_srl3_n_0 ),
        .Q(acc_point_o[10]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1100] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1100]_srl3_n_0 ),
        .Q(acc_point_o[1100]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1101] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1101]_srl3_n_0 ),
        .Q(acc_point_o[1101]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1102] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1102]_srl3_n_0 ),
        .Q(acc_point_o[1102]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1103] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1103]_srl3_n_0 ),
        .Q(acc_point_o[1103]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1104] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1104]_srl3_n_0 ),
        .Q(acc_point_o[1104]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1105] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1105]_srl3_n_0 ),
        .Q(acc_point_o[1105]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1106] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1106]_srl3_n_0 ),
        .Q(acc_point_o[1106]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1107] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1107]_srl3_n_0 ),
        .Q(acc_point_o[1107]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1108] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1108]_srl3_n_0 ),
        .Q(acc_point_o[1108]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1109] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1109]_srl3_n_0 ),
        .Q(acc_point_o[1109]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][110] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][110]_srl3_n_0 ),
        .Q(acc_point_o[110]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1110] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1110]_srl3_n_0 ),
        .Q(acc_point_o[1110]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1111] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1111]_srl3_n_0 ),
        .Q(acc_point_o[1111]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1112] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1112]_srl3_n_0 ),
        .Q(acc_point_o[1112]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1113] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1113]_srl3_n_0 ),
        .Q(acc_point_o[1113]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1114] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1114]_srl3_n_0 ),
        .Q(acc_point_o[1114]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1115] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1115]_srl3_n_0 ),
        .Q(acc_point_o[1115]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1116] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1116]_srl3_n_0 ),
        .Q(acc_point_o[1116]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1117] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1117]_srl3_n_0 ),
        .Q(acc_point_o[1117]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1118] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1118]_srl3_n_0 ),
        .Q(acc_point_o[1118]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1119] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1119]_srl3_n_0 ),
        .Q(acc_point_o[1119]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][111] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][111]_srl3_n_0 ),
        .Q(acc_point_o[111]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1120] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1120]_srl3_n_0 ),
        .Q(acc_point_o[1120]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1121] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1121]_srl3_n_0 ),
        .Q(acc_point_o[1121]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1122] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1122]_srl3_n_0 ),
        .Q(acc_point_o[1122]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1123] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1123]_srl3_n_0 ),
        .Q(acc_point_o[1123]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1124] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1124]_srl3_n_0 ),
        .Q(acc_point_o[1124]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1125] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1125]_srl3_n_0 ),
        .Q(acc_point_o[1125]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1126] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1126]_srl3_n_0 ),
        .Q(acc_point_o[1126]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1127] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1127]_srl3_n_0 ),
        .Q(acc_point_o[1127]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1128] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1128]_srl3_n_0 ),
        .Q(acc_point_o[1128]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1129] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1129]_srl3_n_0 ),
        .Q(acc_point_o[1129]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][112] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][112]_srl3_n_0 ),
        .Q(acc_point_o[112]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1130] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1130]_srl3_n_0 ),
        .Q(acc_point_o[1130]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1131] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1131]_srl3_n_0 ),
        .Q(acc_point_o[1131]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1132] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1132]_srl3_n_0 ),
        .Q(acc_point_o[1132]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1133] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1133]_srl3_n_0 ),
        .Q(acc_point_o[1133]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1134] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1134]_srl3_n_0 ),
        .Q(acc_point_o[1134]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1135] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1135]_srl3_n_0 ),
        .Q(acc_point_o[1135]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1136] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1136]_srl3_n_0 ),
        .Q(acc_point_o[1136]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1137] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1137]_srl3_n_0 ),
        .Q(acc_point_o[1137]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1138] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1138]_srl3_n_0 ),
        .Q(acc_point_o[1138]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1139] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1139]_srl3_n_0 ),
        .Q(acc_point_o[1139]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][113] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][113]_srl3_n_0 ),
        .Q(acc_point_o[113]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1140] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1140]_srl3_n_0 ),
        .Q(acc_point_o[1140]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1141] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1141]_srl3_n_0 ),
        .Q(acc_point_o[1141]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1142] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1142]_srl3_n_0 ),
        .Q(acc_point_o[1142]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1143] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1143]_srl3_n_0 ),
        .Q(acc_point_o[1143]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1144] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1144]_srl3_n_0 ),
        .Q(acc_point_o[1144]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1145] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1145]_srl3_n_0 ),
        .Q(acc_point_o[1145]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1146] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1146]_srl3_n_0 ),
        .Q(acc_point_o[1146]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1147] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1147]_srl3_n_0 ),
        .Q(acc_point_o[1147]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1148] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1148]_srl3_n_0 ),
        .Q(acc_point_o[1148]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1149] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1149]_srl3_n_0 ),
        .Q(acc_point_o[1149]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][114] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][114]_srl3_n_0 ),
        .Q(acc_point_o[114]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1150] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1150]_srl3_n_0 ),
        .Q(acc_point_o[1150]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1151] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1151]_srl3_n_0 ),
        .Q(acc_point_o[1151]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1152] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1152]_srl3_n_0 ),
        .Q(acc_point_o[1152]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1153] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1153]_srl3_n_0 ),
        .Q(acc_point_o[1153]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1154] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1154]_srl3_n_0 ),
        .Q(acc_point_o[1154]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1155] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1155]_srl3_n_0 ),
        .Q(acc_point_o[1155]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1156] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1156]_srl3_n_0 ),
        .Q(acc_point_o[1156]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1157] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1157]_srl3_n_0 ),
        .Q(acc_point_o[1157]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1158] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1158]_srl3_n_0 ),
        .Q(acc_point_o[1158]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1159] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1159]_srl3_n_0 ),
        .Q(acc_point_o[1159]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][115] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][115]_srl3_n_0 ),
        .Q(acc_point_o[115]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1160] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1160]_srl3_n_0 ),
        .Q(acc_point_o[1160]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1161] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1161]_srl3_n_0 ),
        .Q(acc_point_o[1161]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1162] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1162]_srl3_n_0 ),
        .Q(acc_point_o[1162]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1163] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1163]_srl3_n_0 ),
        .Q(acc_point_o[1163]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][116] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][116]_srl3_n_0 ),
        .Q(acc_point_o[116]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][117] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][117]_srl3_n_0 ),
        .Q(acc_point_o[117]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][118] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][118]_srl3_n_0 ),
        .Q(acc_point_o[118]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][119] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][119]_srl3_n_0 ),
        .Q(acc_point_o[119]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][11]_srl3_n_0 ),
        .Q(acc_point_o[11]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][120] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][120]_srl3_n_0 ),
        .Q(acc_point_o[120]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][121] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][121]_srl3_n_0 ),
        .Q(acc_point_o[121]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][122] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][122]_srl3_n_0 ),
        .Q(acc_point_o[122]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][123] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][123]_srl3_n_0 ),
        .Q(acc_point_o[123]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][124] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][124]_srl3_n_0 ),
        .Q(acc_point_o[124]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][125] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][125]_srl3_n_0 ),
        .Q(acc_point_o[125]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][126] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][126]_srl3_n_0 ),
        .Q(acc_point_o[126]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][127] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][127]_srl3_n_0 ),
        .Q(acc_point_o[127]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][128] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][128]_srl3_n_0 ),
        .Q(acc_point_o[128]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][129] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][129]_srl3_n_0 ),
        .Q(acc_point_o[129]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][12]_srl3_n_0 ),
        .Q(acc_point_o[12]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][130] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][130]_srl3_n_0 ),
        .Q(acc_point_o[130]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][131] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][131]_srl3_n_0 ),
        .Q(acc_point_o[131]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][132] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][132]_srl3_n_0 ),
        .Q(acc_point_o[132]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][133] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][133]_srl3_n_0 ),
        .Q(acc_point_o[133]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][134] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][134]_srl3_n_0 ),
        .Q(acc_point_o[134]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][135] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][135]_srl3_n_0 ),
        .Q(acc_point_o[135]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][136] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][136]_srl3_n_0 ),
        .Q(acc_point_o[136]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][137] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][137]_srl3_n_0 ),
        .Q(acc_point_o[137]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][138] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][138]_srl3_n_0 ),
        .Q(acc_point_o[138]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][139] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][139]_srl3_n_0 ),
        .Q(acc_point_o[139]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][13]_srl3_n_0 ),
        .Q(acc_point_o[13]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][140] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][140]_srl3_n_0 ),
        .Q(acc_point_o[140]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][141] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][141]_srl3_n_0 ),
        .Q(acc_point_o[141]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][142] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][142]_srl3_n_0 ),
        .Q(acc_point_o[142]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][143] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][143]_srl3_n_0 ),
        .Q(acc_point_o[143]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][144] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][144]_srl3_n_0 ),
        .Q(acc_point_o[144]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][145] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][145]_srl3_n_0 ),
        .Q(acc_point_o[145]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][146] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][146]_srl3_n_0 ),
        .Q(acc_point_o[146]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][147] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][147]_srl3_n_0 ),
        .Q(acc_point_o[147]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][148] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][148]_srl3_n_0 ),
        .Q(acc_point_o[148]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][149] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][149]_srl3_n_0 ),
        .Q(acc_point_o[149]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][14]_srl3_n_0 ),
        .Q(acc_point_o[14]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][150] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][150]_srl3_n_0 ),
        .Q(acc_point_o[150]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][151] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][151]_srl3_n_0 ),
        .Q(acc_point_o[151]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][152] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][152]_srl3_n_0 ),
        .Q(acc_point_o[152]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][153] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][153]_srl3_n_0 ),
        .Q(acc_point_o[153]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][154] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][154]_srl3_n_0 ),
        .Q(acc_point_o[154]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][155] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][155]_srl3_n_0 ),
        .Q(acc_point_o[155]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][156] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][156]_srl3_n_0 ),
        .Q(acc_point_o[156]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][157] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][157]_srl3_n_0 ),
        .Q(acc_point_o[157]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][158] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][158]_srl3_n_0 ),
        .Q(acc_point_o[158]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][159] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][159]_srl3_n_0 ),
        .Q(acc_point_o[159]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][15]_srl3_n_0 ),
        .Q(acc_point_o[15]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][160] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][160]_srl3_n_0 ),
        .Q(acc_point_o[160]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][161] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][161]_srl3_n_0 ),
        .Q(acc_point_o[161]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][162] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][162]_srl3_n_0 ),
        .Q(acc_point_o[162]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][163] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][163]_srl3_n_0 ),
        .Q(acc_point_o[163]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][164] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][164]_srl3_n_0 ),
        .Q(acc_point_o[164]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][165] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][165]_srl3_n_0 ),
        .Q(acc_point_o[165]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][166] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][166]_srl3_n_0 ),
        .Q(acc_point_o[166]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][167] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][167]_srl3_n_0 ),
        .Q(acc_point_o[167]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][168] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][168]_srl3_n_0 ),
        .Q(acc_point_o[168]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][169] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][169]_srl3_n_0 ),
        .Q(acc_point_o[169]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][16]_srl3_n_0 ),
        .Q(acc_point_o[16]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][170] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][170]_srl3_n_0 ),
        .Q(acc_point_o[170]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][171] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][171]_srl3_n_0 ),
        .Q(acc_point_o[171]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][172] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][172]_srl3_n_0 ),
        .Q(acc_point_o[172]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][173] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][173]_srl3_n_0 ),
        .Q(acc_point_o[173]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][174] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][174]_srl3_n_0 ),
        .Q(acc_point_o[174]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][175] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][175]_srl3_n_0 ),
        .Q(acc_point_o[175]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][176] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][176]_srl3_n_0 ),
        .Q(acc_point_o[176]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][177] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][177]_srl3_n_0 ),
        .Q(acc_point_o[177]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][178] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][178]_srl3_n_0 ),
        .Q(acc_point_o[178]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][179] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][179]_srl3_n_0 ),
        .Q(acc_point_o[179]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][17]_srl3_n_0 ),
        .Q(acc_point_o[17]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][180] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][180]_srl3_n_0 ),
        .Q(acc_point_o[180]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][181] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][181]_srl3_n_0 ),
        .Q(acc_point_o[181]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][182] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][182]_srl3_n_0 ),
        .Q(acc_point_o[182]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][183] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][183]_srl3_n_0 ),
        .Q(acc_point_o[183]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][184] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][184]_srl3_n_0 ),
        .Q(acc_point_o[184]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][185] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][185]_srl3_n_0 ),
        .Q(acc_point_o[185]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][186] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][186]_srl3_n_0 ),
        .Q(acc_point_o[186]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][187] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][187]_srl3_n_0 ),
        .Q(acc_point_o[187]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][188] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][188]_srl3_n_0 ),
        .Q(acc_point_o[188]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][189] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][189]_srl3_n_0 ),
        .Q(acc_point_o[189]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][18]_srl3_n_0 ),
        .Q(acc_point_o[18]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][190] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][190]_srl3_n_0 ),
        .Q(acc_point_o[190]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][191] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][191]_srl3_n_0 ),
        .Q(acc_point_o[191]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][192] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][192]_srl3_n_0 ),
        .Q(acc_point_o[192]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][193] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][193]_srl3_n_0 ),
        .Q(acc_point_o[193]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][194] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][194]_srl3_n_0 ),
        .Q(acc_point_o[194]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][195] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][195]_srl3_n_0 ),
        .Q(acc_point_o[195]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][196] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][196]_srl3_n_0 ),
        .Q(acc_point_o[196]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][197] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][197]_srl3_n_0 ),
        .Q(acc_point_o[197]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][198] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][198]_srl3_n_0 ),
        .Q(acc_point_o[198]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][199] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][199]_srl3_n_0 ),
        .Q(acc_point_o[199]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][19]_srl3_n_0 ),
        .Q(acc_point_o[19]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][1]_srl3_n_0 ),
        .Q(acc_point_o[1]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][200] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][200]_srl3_n_0 ),
        .Q(acc_point_o[200]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][201] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][201]_srl3_n_0 ),
        .Q(acc_point_o[201]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][202] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][202]_srl3_n_0 ),
        .Q(acc_point_o[202]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][203] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][203]_srl3_n_0 ),
        .Q(acc_point_o[203]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][204] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][204]_srl3_n_0 ),
        .Q(acc_point_o[204]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][205] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][205]_srl3_n_0 ),
        .Q(acc_point_o[205]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][206] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][206]_srl3_n_0 ),
        .Q(acc_point_o[206]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][207] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][207]_srl3_n_0 ),
        .Q(acc_point_o[207]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][208] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][208]_srl3_n_0 ),
        .Q(acc_point_o[208]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][209] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][209]_srl3_n_0 ),
        .Q(acc_point_o[209]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][20]_srl3_n_0 ),
        .Q(acc_point_o[20]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][210] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][210]_srl3_n_0 ),
        .Q(acc_point_o[210]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][211] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][211]_srl3_n_0 ),
        .Q(acc_point_o[211]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][212] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][212]_srl3_n_0 ),
        .Q(acc_point_o[212]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][213] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][213]_srl3_n_0 ),
        .Q(acc_point_o[213]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][214] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][214]_srl3_n_0 ),
        .Q(acc_point_o[214]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][215] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][215]_srl3_n_0 ),
        .Q(acc_point_o[215]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][216] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][216]_srl3_n_0 ),
        .Q(acc_point_o[216]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][217] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][217]_srl3_n_0 ),
        .Q(acc_point_o[217]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][218] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][218]_srl3_n_0 ),
        .Q(acc_point_o[218]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][219] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][219]_srl3_n_0 ),
        .Q(acc_point_o[219]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][21]_srl3_n_0 ),
        .Q(acc_point_o[21]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][220] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][220]_srl3_n_0 ),
        .Q(acc_point_o[220]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][221] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][221]_srl3_n_0 ),
        .Q(acc_point_o[221]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][222] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][222]_srl3_n_0 ),
        .Q(acc_point_o[222]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][223] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][223]_srl3_n_0 ),
        .Q(acc_point_o[223]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][224] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][224]_srl3_n_0 ),
        .Q(acc_point_o[224]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][225] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][225]_srl3_n_0 ),
        .Q(acc_point_o[225]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][226] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][226]_srl3_n_0 ),
        .Q(acc_point_o[226]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][227] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][227]_srl3_n_0 ),
        .Q(acc_point_o[227]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][228] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][228]_srl3_n_0 ),
        .Q(acc_point_o[228]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][229] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][229]_srl3_n_0 ),
        .Q(acc_point_o[229]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][22]_srl3_n_0 ),
        .Q(acc_point_o[22]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][230] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][230]_srl3_n_0 ),
        .Q(acc_point_o[230]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][231] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][231]_srl3_n_0 ),
        .Q(acc_point_o[231]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][232] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][232]_srl3_n_0 ),
        .Q(acc_point_o[232]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][233] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][233]_srl3_n_0 ),
        .Q(acc_point_o[233]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][234] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][234]_srl3_n_0 ),
        .Q(acc_point_o[234]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][235] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][235]_srl3_n_0 ),
        .Q(acc_point_o[235]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][236] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][236]_srl3_n_0 ),
        .Q(acc_point_o[236]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][237] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][237]_srl3_n_0 ),
        .Q(acc_point_o[237]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][238] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][238]_srl3_n_0 ),
        .Q(acc_point_o[238]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][239] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][239]_srl3_n_0 ),
        .Q(acc_point_o[239]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][23]_srl3_n_0 ),
        .Q(acc_point_o[23]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][240] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][240]_srl3_n_0 ),
        .Q(acc_point_o[240]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][241] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][241]_srl3_n_0 ),
        .Q(acc_point_o[241]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][242] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][242]_srl3_n_0 ),
        .Q(acc_point_o[242]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][243] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][243]_srl3_n_0 ),
        .Q(acc_point_o[243]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][244] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][244]_srl3_n_0 ),
        .Q(acc_point_o[244]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][245] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][245]_srl3_n_0 ),
        .Q(acc_point_o[245]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][246] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][246]_srl3_n_0 ),
        .Q(acc_point_o[246]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][247] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][247]_srl3_n_0 ),
        .Q(acc_point_o[247]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][248] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][248]_srl3_n_0 ),
        .Q(acc_point_o[248]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][249] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][249]_srl3_n_0 ),
        .Q(acc_point_o[249]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][24]_srl3_n_0 ),
        .Q(acc_point_o[24]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][250] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][250]_srl3_n_0 ),
        .Q(acc_point_o[250]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][251] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][251]_srl3_n_0 ),
        .Q(acc_point_o[251]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][252] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][252]_srl3_n_0 ),
        .Q(acc_point_o[252]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][253] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][253]_srl3_n_0 ),
        .Q(acc_point_o[253]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][254] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][254]_srl3_n_0 ),
        .Q(acc_point_o[254]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][255] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][255]_srl3_n_0 ),
        .Q(acc_point_o[255]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][256] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][256]_srl3_n_0 ),
        .Q(acc_point_o[256]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][257] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][257]_srl3_n_0 ),
        .Q(acc_point_o[257]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][258] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][258]_srl3_n_0 ),
        .Q(acc_point_o[258]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][259] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][259]_srl3_n_0 ),
        .Q(acc_point_o[259]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][25]_srl3_n_0 ),
        .Q(acc_point_o[25]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][260] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][260]_srl3_n_0 ),
        .Q(acc_point_o[260]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][261] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][261]_srl3_n_0 ),
        .Q(acc_point_o[261]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][262] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][262]_srl3_n_0 ),
        .Q(acc_point_o[262]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][263] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][263]_srl3_n_0 ),
        .Q(acc_point_o[263]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][264] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][264]_srl3_n_0 ),
        .Q(acc_point_o[264]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][265] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][265]_srl3_n_0 ),
        .Q(acc_point_o[265]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][266] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][266]_srl3_n_0 ),
        .Q(acc_point_o[266]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][267] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][267]_srl3_n_0 ),
        .Q(acc_point_o[267]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][268] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][268]_srl3_n_0 ),
        .Q(acc_point_o[268]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][269] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][269]_srl3_n_0 ),
        .Q(acc_point_o[269]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][26]_srl3_n_0 ),
        .Q(acc_point_o[26]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][270] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][270]_srl3_n_0 ),
        .Q(acc_point_o[270]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][271] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][271]_srl3_n_0 ),
        .Q(acc_point_o[271]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][272] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][272]_srl3_n_0 ),
        .Q(acc_point_o[272]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][273] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][273]_srl3_n_0 ),
        .Q(acc_point_o[273]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][274] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][274]_srl3_n_0 ),
        .Q(acc_point_o[274]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][275] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][275]_srl3_n_0 ),
        .Q(acc_point_o[275]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][276] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][276]_srl3_n_0 ),
        .Q(acc_point_o[276]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][277] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][277]_srl3_n_0 ),
        .Q(acc_point_o[277]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][278] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][278]_srl3_n_0 ),
        .Q(acc_point_o[278]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][279] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][279]_srl3_n_0 ),
        .Q(acc_point_o[279]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][27]_srl3_n_0 ),
        .Q(acc_point_o[27]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][280] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][280]_srl3_n_0 ),
        .Q(acc_point_o[280]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][281] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][281]_srl3_n_0 ),
        .Q(acc_point_o[281]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][282] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][282]_srl3_n_0 ),
        .Q(acc_point_o[282]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][283] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][283]_srl3_n_0 ),
        .Q(acc_point_o[283]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][284] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][284]_srl3_n_0 ),
        .Q(acc_point_o[284]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][285] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][285]_srl3_n_0 ),
        .Q(acc_point_o[285]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][286] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][286]_srl3_n_0 ),
        .Q(acc_point_o[286]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][287] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][287]_srl3_n_0 ),
        .Q(acc_point_o[287]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][288] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][288]_srl3_n_0 ),
        .Q(acc_point_o[288]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][289] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][289]_srl3_n_0 ),
        .Q(acc_point_o[289]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][28]_srl3_n_0 ),
        .Q(acc_point_o[28]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][290] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][290]_srl3_n_0 ),
        .Q(acc_point_o[290]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][291] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][291]_srl3_n_0 ),
        .Q(acc_point_o[291]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][292] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][292]_srl3_n_0 ),
        .Q(acc_point_o[292]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][293] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][293]_srl3_n_0 ),
        .Q(acc_point_o[293]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][294] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][294]_srl3_n_0 ),
        .Q(acc_point_o[294]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][295] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][295]_srl3_n_0 ),
        .Q(acc_point_o[295]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][296] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][296]_srl3_n_0 ),
        .Q(acc_point_o[296]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][297] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][297]_srl3_n_0 ),
        .Q(acc_point_o[297]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][298] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][298]_srl3_n_0 ),
        .Q(acc_point_o[298]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][299] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][299]_srl3_n_0 ),
        .Q(acc_point_o[299]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][29]_srl3_n_0 ),
        .Q(acc_point_o[29]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][2]_srl3_n_0 ),
        .Q(acc_point_o[2]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][300] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][300]_srl3_n_0 ),
        .Q(acc_point_o[300]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][301] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][301]_srl3_n_0 ),
        .Q(acc_point_o[301]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][302] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][302]_srl3_n_0 ),
        .Q(acc_point_o[302]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][303] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][303]_srl3_n_0 ),
        .Q(acc_point_o[303]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][304] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][304]_srl3_n_0 ),
        .Q(acc_point_o[304]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][305] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][305]_srl3_n_0 ),
        .Q(acc_point_o[305]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][306] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][306]_srl3_n_0 ),
        .Q(acc_point_o[306]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][307] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][307]_srl3_n_0 ),
        .Q(acc_point_o[307]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][308] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][308]_srl3_n_0 ),
        .Q(acc_point_o[308]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][309] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][309]_srl3_n_0 ),
        .Q(acc_point_o[309]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][30]_srl3_n_0 ),
        .Q(acc_point_o[30]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][310] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][310]_srl3_n_0 ),
        .Q(acc_point_o[310]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][311] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][311]_srl3_n_0 ),
        .Q(acc_point_o[311]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][312] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][312]_srl3_n_0 ),
        .Q(acc_point_o[312]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][313] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][313]_srl3_n_0 ),
        .Q(acc_point_o[313]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][314] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][314]_srl3_n_0 ),
        .Q(acc_point_o[314]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][315] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][315]_srl3_n_0 ),
        .Q(acc_point_o[315]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][316] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][316]_srl3_n_0 ),
        .Q(acc_point_o[316]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][317] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][317]_srl3_n_0 ),
        .Q(acc_point_o[317]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][318] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][318]_srl3_n_0 ),
        .Q(acc_point_o[318]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][319] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][319]_srl3_n_0 ),
        .Q(acc_point_o[319]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][31]_srl3_n_0 ),
        .Q(acc_point_o[31]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][320] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][320]_srl3_n_0 ),
        .Q(acc_point_o[320]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][321] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][321]_srl3_n_0 ),
        .Q(acc_point_o[321]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][322] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][322]_srl3_n_0 ),
        .Q(acc_point_o[322]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][323] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][323]_srl3_n_0 ),
        .Q(acc_point_o[323]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][324] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][324]_srl3_n_0 ),
        .Q(acc_point_o[324]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][325] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][325]_srl3_n_0 ),
        .Q(acc_point_o[325]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][326] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][326]_srl3_n_0 ),
        .Q(acc_point_o[326]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][327] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][327]_srl3_n_0 ),
        .Q(acc_point_o[327]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][328] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][328]_srl3_n_0 ),
        .Q(acc_point_o[328]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][329] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][329]_srl3_n_0 ),
        .Q(acc_point_o[329]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][32] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][32]_srl3_n_0 ),
        .Q(acc_point_o[32]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][330] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][330]_srl3_n_0 ),
        .Q(acc_point_o[330]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][331] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][331]_srl3_n_0 ),
        .Q(acc_point_o[331]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][332] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][332]_srl3_n_0 ),
        .Q(acc_point_o[332]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][333] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][333]_srl3_n_0 ),
        .Q(acc_point_o[333]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][334] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][334]_srl3_n_0 ),
        .Q(acc_point_o[334]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][335] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][335]_srl3_n_0 ),
        .Q(acc_point_o[335]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][336] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][336]_srl3_n_0 ),
        .Q(acc_point_o[336]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][337] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][337]_srl3_n_0 ),
        .Q(acc_point_o[337]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][338] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][338]_srl3_n_0 ),
        .Q(acc_point_o[338]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][339] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][339]_srl3_n_0 ),
        .Q(acc_point_o[339]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][33] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][33]_srl3_n_0 ),
        .Q(acc_point_o[33]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][340] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][340]_srl3_n_0 ),
        .Q(acc_point_o[340]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][341] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][341]_srl3_n_0 ),
        .Q(acc_point_o[341]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][342] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][342]_srl3_n_0 ),
        .Q(acc_point_o[342]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][343] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][343]_srl3_n_0 ),
        .Q(acc_point_o[343]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][344] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][344]_srl3_n_0 ),
        .Q(acc_point_o[344]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][345] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][345]_srl3_n_0 ),
        .Q(acc_point_o[345]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][346] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][346]_srl3_n_0 ),
        .Q(acc_point_o[346]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][347] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][347]_srl3_n_0 ),
        .Q(acc_point_o[347]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][348] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][348]_srl3_n_0 ),
        .Q(acc_point_o[348]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][349] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][349]_srl3_n_0 ),
        .Q(acc_point_o[349]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][34] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][34]_srl3_n_0 ),
        .Q(acc_point_o[34]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][350] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][350]_srl3_n_0 ),
        .Q(acc_point_o[350]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][351] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][351]_srl3_n_0 ),
        .Q(acc_point_o[351]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][352] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][352]_srl3_n_0 ),
        .Q(acc_point_o[352]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][353] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][353]_srl3_n_0 ),
        .Q(acc_point_o[353]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][354] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][354]_srl3_n_0 ),
        .Q(acc_point_o[354]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][355] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][355]_srl3_n_0 ),
        .Q(acc_point_o[355]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][356] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][356]_srl3_n_0 ),
        .Q(acc_point_o[356]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][357] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][357]_srl3_n_0 ),
        .Q(acc_point_o[357]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][358] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][358]_srl3_n_0 ),
        .Q(acc_point_o[358]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][359] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][359]_srl3_n_0 ),
        .Q(acc_point_o[359]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][35] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][35]_srl3_n_0 ),
        .Q(acc_point_o[35]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][360] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][360]_srl3_n_0 ),
        .Q(acc_point_o[360]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][361] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][361]_srl3_n_0 ),
        .Q(acc_point_o[361]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][362] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][362]_srl3_n_0 ),
        .Q(acc_point_o[362]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][363] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][363]_srl3_n_0 ),
        .Q(acc_point_o[363]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][364] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][364]_srl3_n_0 ),
        .Q(acc_point_o[364]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][365] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][365]_srl3_n_0 ),
        .Q(acc_point_o[365]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][366] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][366]_srl3_n_0 ),
        .Q(acc_point_o[366]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][367] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][367]_srl3_n_0 ),
        .Q(acc_point_o[367]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][368] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][368]_srl3_n_0 ),
        .Q(acc_point_o[368]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][369] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][369]_srl3_n_0 ),
        .Q(acc_point_o[369]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][36] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][36]_srl3_n_0 ),
        .Q(acc_point_o[36]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][370] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][370]_srl3_n_0 ),
        .Q(acc_point_o[370]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][371] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][371]_srl3_n_0 ),
        .Q(acc_point_o[371]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][372] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][372]_srl3_n_0 ),
        .Q(acc_point_o[372]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][373] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][373]_srl3_n_0 ),
        .Q(acc_point_o[373]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][374] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][374]_srl3_n_0 ),
        .Q(acc_point_o[374]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][375] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][375]_srl3_n_0 ),
        .Q(acc_point_o[375]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][376] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][376]_srl3_n_0 ),
        .Q(acc_point_o[376]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][377] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][377]_srl3_n_0 ),
        .Q(acc_point_o[377]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][378] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][378]_srl3_n_0 ),
        .Q(acc_point_o[378]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][379] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][379]_srl3_n_0 ),
        .Q(acc_point_o[379]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][37] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][37]_srl3_n_0 ),
        .Q(acc_point_o[37]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][380] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][380]_srl3_n_0 ),
        .Q(acc_point_o[380]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][381] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][381]_srl3_n_0 ),
        .Q(acc_point_o[381]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][382] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][382]_srl3_n_0 ),
        .Q(acc_point_o[382]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][383] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][383]_srl3_n_0 ),
        .Q(acc_point_o[383]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][384] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][384]_srl3_n_0 ),
        .Q(acc_point_o[384]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][385] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][385]_srl3_n_0 ),
        .Q(acc_point_o[385]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][386] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][386]_srl3_n_0 ),
        .Q(acc_point_o[386]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][387] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][387]_srl3_n_0 ),
        .Q(acc_point_o[387]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][388] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][388]_srl3_n_0 ),
        .Q(acc_point_o[388]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][389] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][389]_srl3_n_0 ),
        .Q(acc_point_o[389]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][38] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][38]_srl3_n_0 ),
        .Q(acc_point_o[38]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][390] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][390]_srl3_n_0 ),
        .Q(acc_point_o[390]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][391] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][391]_srl3_n_0 ),
        .Q(acc_point_o[391]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][392] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][392]_srl3_n_0 ),
        .Q(acc_point_o[392]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][393] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][393]_srl3_n_0 ),
        .Q(acc_point_o[393]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][394] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][394]_srl3_n_0 ),
        .Q(acc_point_o[394]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][395] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][395]_srl3_n_0 ),
        .Q(acc_point_o[395]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][396] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][396]_srl3_n_0 ),
        .Q(acc_point_o[396]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][397] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][397]_srl3_n_0 ),
        .Q(acc_point_o[397]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][398] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][398]_srl3_n_0 ),
        .Q(acc_point_o[398]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][399] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][399]_srl3_n_0 ),
        .Q(acc_point_o[399]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][39] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][39]_srl3_n_0 ),
        .Q(acc_point_o[39]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][3]_srl3_n_0 ),
        .Q(acc_point_o[3]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][400] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][400]_srl3_n_0 ),
        .Q(acc_point_o[400]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][401] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][401]_srl3_n_0 ),
        .Q(acc_point_o[401]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][402] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][402]_srl3_n_0 ),
        .Q(acc_point_o[402]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][403] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][403]_srl3_n_0 ),
        .Q(acc_point_o[403]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][404] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][404]_srl3_n_0 ),
        .Q(acc_point_o[404]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][405] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][405]_srl3_n_0 ),
        .Q(acc_point_o[405]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][406] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][406]_srl3_n_0 ),
        .Q(acc_point_o[406]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][407] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][407]_srl3_n_0 ),
        .Q(acc_point_o[407]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][408] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][408]_srl3_n_0 ),
        .Q(acc_point_o[408]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][409] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][409]_srl3_n_0 ),
        .Q(acc_point_o[409]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][40] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][40]_srl3_n_0 ),
        .Q(acc_point_o[40]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][410] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][410]_srl3_n_0 ),
        .Q(acc_point_o[410]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][411] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][411]_srl3_n_0 ),
        .Q(acc_point_o[411]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][412] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][412]_srl3_n_0 ),
        .Q(acc_point_o[412]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][413] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][413]_srl3_n_0 ),
        .Q(acc_point_o[413]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][414] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][414]_srl3_n_0 ),
        .Q(acc_point_o[414]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][415] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][415]_srl3_n_0 ),
        .Q(acc_point_o[415]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][416] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][416]_srl3_n_0 ),
        .Q(acc_point_o[416]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][417] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][417]_srl3_n_0 ),
        .Q(acc_point_o[417]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][418] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][418]_srl3_n_0 ),
        .Q(acc_point_o[418]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][419] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][419]_srl3_n_0 ),
        .Q(acc_point_o[419]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][41] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][41]_srl3_n_0 ),
        .Q(acc_point_o[41]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][420] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][420]_srl3_n_0 ),
        .Q(acc_point_o[420]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][421] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][421]_srl3_n_0 ),
        .Q(acc_point_o[421]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][422] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][422]_srl3_n_0 ),
        .Q(acc_point_o[422]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][423] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][423]_srl3_n_0 ),
        .Q(acc_point_o[423]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][424] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][424]_srl3_n_0 ),
        .Q(acc_point_o[424]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][425] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][425]_srl3_n_0 ),
        .Q(acc_point_o[425]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][426] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][426]_srl3_n_0 ),
        .Q(acc_point_o[426]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][427] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][427]_srl3_n_0 ),
        .Q(acc_point_o[427]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][428] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][428]_srl3_n_0 ),
        .Q(acc_point_o[428]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][429] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][429]_srl3_n_0 ),
        .Q(acc_point_o[429]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][42] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][42]_srl3_n_0 ),
        .Q(acc_point_o[42]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][430] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][430]_srl3_n_0 ),
        .Q(acc_point_o[430]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][431] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][431]_srl3_n_0 ),
        .Q(acc_point_o[431]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][432] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][432]_srl3_n_0 ),
        .Q(acc_point_o[432]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][433] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][433]_srl3_n_0 ),
        .Q(acc_point_o[433]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][434] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][434]_srl3_n_0 ),
        .Q(acc_point_o[434]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][435] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][435]_srl3_n_0 ),
        .Q(acc_point_o[435]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][436] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][436]_srl3_n_0 ),
        .Q(acc_point_o[436]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][437] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][437]_srl3_n_0 ),
        .Q(acc_point_o[437]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][438] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][438]_srl3_n_0 ),
        .Q(acc_point_o[438]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][439] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][439]_srl3_n_0 ),
        .Q(acc_point_o[439]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][43] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][43]_srl3_n_0 ),
        .Q(acc_point_o[43]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][440] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][440]_srl3_n_0 ),
        .Q(acc_point_o[440]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][441] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][441]_srl3_n_0 ),
        .Q(acc_point_o[441]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][442] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][442]_srl3_n_0 ),
        .Q(acc_point_o[442]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][443] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][443]_srl3_n_0 ),
        .Q(acc_point_o[443]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][444] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][444]_srl3_n_0 ),
        .Q(acc_point_o[444]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][445] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][445]_srl3_n_0 ),
        .Q(acc_point_o[445]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][446] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][446]_srl3_n_0 ),
        .Q(acc_point_o[446]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][447] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][447]_srl3_n_0 ),
        .Q(acc_point_o[447]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][448] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][448]_srl3_n_0 ),
        .Q(acc_point_o[448]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][449] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][449]_srl3_n_0 ),
        .Q(acc_point_o[449]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][44] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][44]_srl3_n_0 ),
        .Q(acc_point_o[44]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][450] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][450]_srl3_n_0 ),
        .Q(acc_point_o[450]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][451] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][451]_srl3_n_0 ),
        .Q(acc_point_o[451]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][452] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][452]_srl3_n_0 ),
        .Q(acc_point_o[452]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][453] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][453]_srl3_n_0 ),
        .Q(acc_point_o[453]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][454] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][454]_srl3_n_0 ),
        .Q(acc_point_o[454]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][455] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][455]_srl3_n_0 ),
        .Q(acc_point_o[455]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][456] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][456]_srl3_n_0 ),
        .Q(acc_point_o[456]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][457] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][457]_srl3_n_0 ),
        .Q(acc_point_o[457]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][458] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][458]_srl3_n_0 ),
        .Q(acc_point_o[458]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][459] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][459]_srl3_n_0 ),
        .Q(acc_point_o[459]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][45] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][45]_srl3_n_0 ),
        .Q(acc_point_o[45]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][460] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][460]_srl3_n_0 ),
        .Q(acc_point_o[460]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][461] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][461]_srl3_n_0 ),
        .Q(acc_point_o[461]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][462] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][462]_srl3_n_0 ),
        .Q(acc_point_o[462]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][463] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][463]_srl3_n_0 ),
        .Q(acc_point_o[463]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][464] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][464]_srl3_n_0 ),
        .Q(acc_point_o[464]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][465] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][465]_srl3_n_0 ),
        .Q(acc_point_o[465]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][466] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][466]_srl3_n_0 ),
        .Q(acc_point_o[466]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][467] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][467]_srl3_n_0 ),
        .Q(acc_point_o[467]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][468] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][468]_srl3_n_0 ),
        .Q(acc_point_o[468]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][469] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][469]_srl3_n_0 ),
        .Q(acc_point_o[469]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][46] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][46]_srl3_n_0 ),
        .Q(acc_point_o[46]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][470] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][470]_srl3_n_0 ),
        .Q(acc_point_o[470]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][471] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][471]_srl3_n_0 ),
        .Q(acc_point_o[471]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][472] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][472]_srl3_n_0 ),
        .Q(acc_point_o[472]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][473] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][473]_srl3_n_0 ),
        .Q(acc_point_o[473]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][474] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][474]_srl3_n_0 ),
        .Q(acc_point_o[474]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][475] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][475]_srl3_n_0 ),
        .Q(acc_point_o[475]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][476] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][476]_srl3_n_0 ),
        .Q(acc_point_o[476]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][477] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][477]_srl3_n_0 ),
        .Q(acc_point_o[477]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][478] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][478]_srl3_n_0 ),
        .Q(acc_point_o[478]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][479] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][479]_srl3_n_0 ),
        .Q(acc_point_o[479]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][47] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][47]_srl3_n_0 ),
        .Q(acc_point_o[47]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][480] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][480]_srl3_n_0 ),
        .Q(acc_point_o[480]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][481] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][481]_srl3_n_0 ),
        .Q(acc_point_o[481]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][482] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][482]_srl3_n_0 ),
        .Q(acc_point_o[482]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][483] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][483]_srl3_n_0 ),
        .Q(acc_point_o[483]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][484] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][484]_srl3_n_0 ),
        .Q(acc_point_o[484]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][485] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][485]_srl3_n_0 ),
        .Q(acc_point_o[485]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][486] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][486]_srl3_n_0 ),
        .Q(acc_point_o[486]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][487] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][487]_srl3_n_0 ),
        .Q(acc_point_o[487]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][488] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][488]_srl3_n_0 ),
        .Q(acc_point_o[488]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][489] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][489]_srl3_n_0 ),
        .Q(acc_point_o[489]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][48] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][48]_srl3_n_0 ),
        .Q(acc_point_o[48]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][490] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][490]_srl3_n_0 ),
        .Q(acc_point_o[490]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][491] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][491]_srl3_n_0 ),
        .Q(acc_point_o[491]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][492] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][492]_srl3_n_0 ),
        .Q(acc_point_o[492]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][493] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][493]_srl3_n_0 ),
        .Q(acc_point_o[493]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][494] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][494]_srl3_n_0 ),
        .Q(acc_point_o[494]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][495] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][495]_srl3_n_0 ),
        .Q(acc_point_o[495]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][496] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][496]_srl3_n_0 ),
        .Q(acc_point_o[496]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][497] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][497]_srl3_n_0 ),
        .Q(acc_point_o[497]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][498] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][498]_srl3_n_0 ),
        .Q(acc_point_o[498]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][499] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][499]_srl3_n_0 ),
        .Q(acc_point_o[499]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][49] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][49]_srl3_n_0 ),
        .Q(acc_point_o[49]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][4]_srl3_n_0 ),
        .Q(acc_point_o[4]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][500] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][500]_srl3_n_0 ),
        .Q(acc_point_o[500]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][501] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][501]_srl3_n_0 ),
        .Q(acc_point_o[501]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][502] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][502]_srl3_n_0 ),
        .Q(acc_point_o[502]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][503] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][503]_srl3_n_0 ),
        .Q(acc_point_o[503]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][504] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][504]_srl3_n_0 ),
        .Q(acc_point_o[504]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][505] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][505]_srl3_n_0 ),
        .Q(acc_point_o[505]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][506] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][506]_srl3_n_0 ),
        .Q(acc_point_o[506]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][507] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][507]_srl3_n_0 ),
        .Q(acc_point_o[507]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][508] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][508]_srl3_n_0 ),
        .Q(acc_point_o[508]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][509] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][509]_srl3_n_0 ),
        .Q(acc_point_o[509]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][50] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][50]_srl3_n_0 ),
        .Q(acc_point_o[50]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][510] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][510]_srl3_n_0 ),
        .Q(acc_point_o[510]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][511] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][511]_srl3_n_0 ),
        .Q(acc_point_o[511]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][512] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][512]_srl3_n_0 ),
        .Q(acc_point_o[512]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][513] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][513]_srl3_n_0 ),
        .Q(acc_point_o[513]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][514] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][514]_srl3_n_0 ),
        .Q(acc_point_o[514]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][515] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][515]_srl3_n_0 ),
        .Q(acc_point_o[515]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][516] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][516]_srl3_n_0 ),
        .Q(acc_point_o[516]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][517] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][517]_srl3_n_0 ),
        .Q(acc_point_o[517]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][518] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][518]_srl3_n_0 ),
        .Q(acc_point_o[518]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][519] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][519]_srl3_n_0 ),
        .Q(acc_point_o[519]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][51] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][51]_srl3_n_0 ),
        .Q(acc_point_o[51]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][520] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][520]_srl3_n_0 ),
        .Q(acc_point_o[520]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][521] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][521]_srl3_n_0 ),
        .Q(acc_point_o[521]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][522] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][522]_srl3_n_0 ),
        .Q(acc_point_o[522]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][523] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][523]_srl3_n_0 ),
        .Q(acc_point_o[523]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][524] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][524]_srl3_n_0 ),
        .Q(acc_point_o[524]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][525] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][525]_srl3_n_0 ),
        .Q(acc_point_o[525]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][526] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][526]_srl3_n_0 ),
        .Q(acc_point_o[526]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][527] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][527]_srl3_n_0 ),
        .Q(acc_point_o[527]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][528] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][528]_srl3_n_0 ),
        .Q(acc_point_o[528]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][529] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][529]_srl3_n_0 ),
        .Q(acc_point_o[529]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][52] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][52]_srl3_n_0 ),
        .Q(acc_point_o[52]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][530] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][530]_srl3_n_0 ),
        .Q(acc_point_o[530]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][531] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][531]_srl3_n_0 ),
        .Q(acc_point_o[531]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][532] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][532]_srl3_n_0 ),
        .Q(acc_point_o[532]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][533] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][533]_srl3_n_0 ),
        .Q(acc_point_o[533]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][534] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][534]_srl3_n_0 ),
        .Q(acc_point_o[534]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][535] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][535]_srl3_n_0 ),
        .Q(acc_point_o[535]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][536] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][536]_srl3_n_0 ),
        .Q(acc_point_o[536]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][537] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][537]_srl3_n_0 ),
        .Q(acc_point_o[537]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][538] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][538]_srl3_n_0 ),
        .Q(acc_point_o[538]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][539] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][539]_srl3_n_0 ),
        .Q(acc_point_o[539]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][53] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][53]_srl3_n_0 ),
        .Q(acc_point_o[53]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][540] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][540]_srl3_n_0 ),
        .Q(acc_point_o[540]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][541] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][541]_srl3_n_0 ),
        .Q(acc_point_o[541]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][542] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][542]_srl3_n_0 ),
        .Q(acc_point_o[542]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][543] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][543]_srl3_n_0 ),
        .Q(acc_point_o[543]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][544] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][544]_srl3_n_0 ),
        .Q(acc_point_o[544]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][545] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][545]_srl3_n_0 ),
        .Q(acc_point_o[545]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][546] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][546]_srl3_n_0 ),
        .Q(acc_point_o[546]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][547] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][547]_srl3_n_0 ),
        .Q(acc_point_o[547]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][548] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][548]_srl3_n_0 ),
        .Q(acc_point_o[548]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][549] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][549]_srl3_n_0 ),
        .Q(acc_point_o[549]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][54] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][54]_srl3_n_0 ),
        .Q(acc_point_o[54]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][550] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][550]_srl3_n_0 ),
        .Q(acc_point_o[550]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][551] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][551]_srl3_n_0 ),
        .Q(acc_point_o[551]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][552] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][552]_srl3_n_0 ),
        .Q(acc_point_o[552]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][553] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][553]_srl3_n_0 ),
        .Q(acc_point_o[553]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][554] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][554]_srl3_n_0 ),
        .Q(acc_point_o[554]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][555] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][555]_srl3_n_0 ),
        .Q(acc_point_o[555]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][556] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][556]_srl3_n_0 ),
        .Q(acc_point_o[556]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][557] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][557]_srl3_n_0 ),
        .Q(acc_point_o[557]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][558] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][558]_srl3_n_0 ),
        .Q(acc_point_o[558]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][559] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][559]_srl3_n_0 ),
        .Q(acc_point_o[559]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][55] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][55]_srl3_n_0 ),
        .Q(acc_point_o[55]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][560] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][560]_srl3_n_0 ),
        .Q(acc_point_o[560]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][561] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][561]_srl3_n_0 ),
        .Q(acc_point_o[561]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][562] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][562]_srl3_n_0 ),
        .Q(acc_point_o[562]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][563] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][563]_srl3_n_0 ),
        .Q(acc_point_o[563]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][564] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][564]_srl3_n_0 ),
        .Q(acc_point_o[564]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][565] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][565]_srl3_n_0 ),
        .Q(acc_point_o[565]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][566] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][566]_srl3_n_0 ),
        .Q(acc_point_o[566]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][567] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][567]_srl3_n_0 ),
        .Q(acc_point_o[567]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][568] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][568]_srl3_n_0 ),
        .Q(acc_point_o[568]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][569] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][569]_srl3_n_0 ),
        .Q(acc_point_o[569]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][56] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][56]_srl3_n_0 ),
        .Q(acc_point_o[56]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][570] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][570]_srl3_n_0 ),
        .Q(acc_point_o[570]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][571] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][571]_srl3_n_0 ),
        .Q(acc_point_o[571]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][572] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][572]_srl3_n_0 ),
        .Q(acc_point_o[572]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][573] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][573]_srl3_n_0 ),
        .Q(acc_point_o[573]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][574] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][574]_srl3_n_0 ),
        .Q(acc_point_o[574]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][575] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][575]_srl3_n_0 ),
        .Q(acc_point_o[575]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][576] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][576]_srl3_n_0 ),
        .Q(acc_point_o[576]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][577] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][577]_srl3_n_0 ),
        .Q(acc_point_o[577]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][578] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][578]_srl3_n_0 ),
        .Q(acc_point_o[578]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][579] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][579]_srl3_n_0 ),
        .Q(acc_point_o[579]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][57] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][57]_srl3_n_0 ),
        .Q(acc_point_o[57]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][580] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][580]_srl3_n_0 ),
        .Q(acc_point_o[580]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][581] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][581]_srl3_n_0 ),
        .Q(acc_point_o[581]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][582] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][582]_srl3_n_0 ),
        .Q(acc_point_o[582]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][583] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][583]_srl3_n_0 ),
        .Q(acc_point_o[583]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][584] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][584]_srl3_n_0 ),
        .Q(acc_point_o[584]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][585] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][585]_srl3_n_0 ),
        .Q(acc_point_o[585]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][586] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][586]_srl3_n_0 ),
        .Q(acc_point_o[586]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][587] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][587]_srl3_n_0 ),
        .Q(acc_point_o[587]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][588] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][588]_srl3_n_0 ),
        .Q(acc_point_o[588]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][589] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][589]_srl3_n_0 ),
        .Q(acc_point_o[589]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][58] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][58]_srl3_n_0 ),
        .Q(acc_point_o[58]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][590] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][590]_srl3_n_0 ),
        .Q(acc_point_o[590]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][591] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][591]_srl3_n_0 ),
        .Q(acc_point_o[591]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][592] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][592]_srl3_n_0 ),
        .Q(acc_point_o[592]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][593] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][593]_srl3_n_0 ),
        .Q(acc_point_o[593]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][594] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][594]_srl3_n_0 ),
        .Q(acc_point_o[594]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][595] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][595]_srl3_n_0 ),
        .Q(acc_point_o[595]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][596] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][596]_srl3_n_0 ),
        .Q(acc_point_o[596]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][597] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][597]_srl3_n_0 ),
        .Q(acc_point_o[597]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][598] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][598]_srl3_n_0 ),
        .Q(acc_point_o[598]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][599] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][599]_srl3_n_0 ),
        .Q(acc_point_o[599]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][59] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][59]_srl3_n_0 ),
        .Q(acc_point_o[59]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][5]_srl3_n_0 ),
        .Q(acc_point_o[5]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][600] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][600]_srl3_n_0 ),
        .Q(acc_point_o[600]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][601] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][601]_srl3_n_0 ),
        .Q(acc_point_o[601]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][602] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][602]_srl3_n_0 ),
        .Q(acc_point_o[602]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][603] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][603]_srl3_n_0 ),
        .Q(acc_point_o[603]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][604] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][604]_srl3_n_0 ),
        .Q(acc_point_o[604]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][605] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][605]_srl3_n_0 ),
        .Q(acc_point_o[605]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][606] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][606]_srl3_n_0 ),
        .Q(acc_point_o[606]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][607] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][607]_srl3_n_0 ),
        .Q(acc_point_o[607]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][608] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][608]_srl3_n_0 ),
        .Q(acc_point_o[608]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][609] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][609]_srl3_n_0 ),
        .Q(acc_point_o[609]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][60] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][60]_srl3_n_0 ),
        .Q(acc_point_o[60]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][610] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][610]_srl3_n_0 ),
        .Q(acc_point_o[610]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][611] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][611]_srl3_n_0 ),
        .Q(acc_point_o[611]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][612] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][612]_srl3_n_0 ),
        .Q(acc_point_o[612]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][613] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][613]_srl3_n_0 ),
        .Q(acc_point_o[613]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][614] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][614]_srl3_n_0 ),
        .Q(acc_point_o[614]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][615] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][615]_srl3_n_0 ),
        .Q(acc_point_o[615]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][616] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][616]_srl3_n_0 ),
        .Q(acc_point_o[616]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][617] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][617]_srl3_n_0 ),
        .Q(acc_point_o[617]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][618] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][618]_srl3_n_0 ),
        .Q(acc_point_o[618]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][619] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][619]_srl3_n_0 ),
        .Q(acc_point_o[619]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][61] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][61]_srl3_n_0 ),
        .Q(acc_point_o[61]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][620] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][620]_srl3_n_0 ),
        .Q(acc_point_o[620]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][621] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][621]_srl3_n_0 ),
        .Q(acc_point_o[621]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][622] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][622]_srl3_n_0 ),
        .Q(acc_point_o[622]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][623] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][623]_srl3_n_0 ),
        .Q(acc_point_o[623]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][624] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][624]_srl3_n_0 ),
        .Q(acc_point_o[624]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][625] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][625]_srl3_n_0 ),
        .Q(acc_point_o[625]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][626] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][626]_srl3_n_0 ),
        .Q(acc_point_o[626]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][627] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][627]_srl3_n_0 ),
        .Q(acc_point_o[627]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][628] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][628]_srl3_n_0 ),
        .Q(acc_point_o[628]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][629] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][629]_srl3_n_0 ),
        .Q(acc_point_o[629]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][62] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][62]_srl3_n_0 ),
        .Q(acc_point_o[62]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][630] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][630]_srl3_n_0 ),
        .Q(acc_point_o[630]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][631] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][631]_srl3_n_0 ),
        .Q(acc_point_o[631]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][632] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][632]_srl3_n_0 ),
        .Q(acc_point_o[632]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][633] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][633]_srl3_n_0 ),
        .Q(acc_point_o[633]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][634] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][634]_srl3_n_0 ),
        .Q(acc_point_o[634]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][635] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][635]_srl3_n_0 ),
        .Q(acc_point_o[635]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][636] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][636]_srl3_n_0 ),
        .Q(acc_point_o[636]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][637] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][637]_srl3_n_0 ),
        .Q(acc_point_o[637]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][638] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][638]_srl3_n_0 ),
        .Q(acc_point_o[638]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][639] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][639]_srl3_n_0 ),
        .Q(acc_point_o[639]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][63] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][63]_srl3_n_0 ),
        .Q(acc_point_o[63]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][640] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][640]_srl3_n_0 ),
        .Q(acc_point_o[640]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][641] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][641]_srl3_n_0 ),
        .Q(acc_point_o[641]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][642] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][642]_srl3_n_0 ),
        .Q(acc_point_o[642]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][643] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][643]_srl3_n_0 ),
        .Q(acc_point_o[643]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][644] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][644]_srl3_n_0 ),
        .Q(acc_point_o[644]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][645] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][645]_srl3_n_0 ),
        .Q(acc_point_o[645]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][646] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][646]_srl3_n_0 ),
        .Q(acc_point_o[646]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][647] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][647]_srl3_n_0 ),
        .Q(acc_point_o[647]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][648] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][648]_srl3_n_0 ),
        .Q(acc_point_o[648]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][649] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][649]_srl3_n_0 ),
        .Q(acc_point_o[649]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][64] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][64]_srl3_n_0 ),
        .Q(acc_point_o[64]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][650] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][650]_srl3_n_0 ),
        .Q(acc_point_o[650]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][651] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][651]_srl3_n_0 ),
        .Q(acc_point_o[651]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][652] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][652]_srl3_n_0 ),
        .Q(acc_point_o[652]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][653] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][653]_srl3_n_0 ),
        .Q(acc_point_o[653]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][654] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][654]_srl3_n_0 ),
        .Q(acc_point_o[654]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][655] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][655]_srl3_n_0 ),
        .Q(acc_point_o[655]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][656] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][656]_srl3_n_0 ),
        .Q(acc_point_o[656]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][657] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][657]_srl3_n_0 ),
        .Q(acc_point_o[657]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][658] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][658]_srl3_n_0 ),
        .Q(acc_point_o[658]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][659] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][659]_srl3_n_0 ),
        .Q(acc_point_o[659]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][65] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][65]_srl3_n_0 ),
        .Q(acc_point_o[65]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][660] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][660]_srl3_n_0 ),
        .Q(acc_point_o[660]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][661] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][661]_srl3_n_0 ),
        .Q(acc_point_o[661]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][662] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][662]_srl3_n_0 ),
        .Q(acc_point_o[662]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][663] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][663]_srl3_n_0 ),
        .Q(acc_point_o[663]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][664] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][664]_srl3_n_0 ),
        .Q(acc_point_o[664]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][665] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][665]_srl3_n_0 ),
        .Q(acc_point_o[665]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][666] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][666]_srl3_n_0 ),
        .Q(acc_point_o[666]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][667] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][667]_srl3_n_0 ),
        .Q(acc_point_o[667]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][668] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][668]_srl3_n_0 ),
        .Q(acc_point_o[668]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][669] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][669]_srl3_n_0 ),
        .Q(acc_point_o[669]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][66] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][66]_srl3_n_0 ),
        .Q(acc_point_o[66]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][670] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][670]_srl3_n_0 ),
        .Q(acc_point_o[670]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][671] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][671]_srl3_n_0 ),
        .Q(acc_point_o[671]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][672] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][672]_srl3_n_0 ),
        .Q(acc_point_o[672]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][673] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][673]_srl3_n_0 ),
        .Q(acc_point_o[673]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][674] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][674]_srl3_n_0 ),
        .Q(acc_point_o[674]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][675] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][675]_srl3_n_0 ),
        .Q(acc_point_o[675]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][676] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][676]_srl3_n_0 ),
        .Q(acc_point_o[676]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][677] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][677]_srl3_n_0 ),
        .Q(acc_point_o[677]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][678] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][678]_srl3_n_0 ),
        .Q(acc_point_o[678]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][679] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][679]_srl3_n_0 ),
        .Q(acc_point_o[679]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][67] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][67]_srl3_n_0 ),
        .Q(acc_point_o[67]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][680] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][680]_srl3_n_0 ),
        .Q(acc_point_o[680]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][681] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][681]_srl3_n_0 ),
        .Q(acc_point_o[681]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][682] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][682]_srl3_n_0 ),
        .Q(acc_point_o[682]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][683] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][683]_srl3_n_0 ),
        .Q(acc_point_o[683]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][684] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][684]_srl3_n_0 ),
        .Q(acc_point_o[684]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][685] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][685]_srl3_n_0 ),
        .Q(acc_point_o[685]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][686] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][686]_srl3_n_0 ),
        .Q(acc_point_o[686]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][687] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][687]_srl3_n_0 ),
        .Q(acc_point_o[687]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][688] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][688]_srl3_n_0 ),
        .Q(acc_point_o[688]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][689] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][689]_srl3_n_0 ),
        .Q(acc_point_o[689]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][68] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][68]_srl3_n_0 ),
        .Q(acc_point_o[68]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][690] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][690]_srl3_n_0 ),
        .Q(acc_point_o[690]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][691] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][691]_srl3_n_0 ),
        .Q(acc_point_o[691]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][692] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][692]_srl3_n_0 ),
        .Q(acc_point_o[692]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][693] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][693]_srl3_n_0 ),
        .Q(acc_point_o[693]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][694] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][694]_srl3_n_0 ),
        .Q(acc_point_o[694]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][695] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][695]_srl3_n_0 ),
        .Q(acc_point_o[695]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][696] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][696]_srl3_n_0 ),
        .Q(acc_point_o[696]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][697] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][697]_srl3_n_0 ),
        .Q(acc_point_o[697]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][698] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][698]_srl3_n_0 ),
        .Q(acc_point_o[698]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][699] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][699]_srl3_n_0 ),
        .Q(acc_point_o[699]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][69] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][69]_srl3_n_0 ),
        .Q(acc_point_o[69]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][6]_srl3_n_0 ),
        .Q(acc_point_o[6]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][700] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][700]_srl3_n_0 ),
        .Q(acc_point_o[700]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][701] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][701]_srl3_n_0 ),
        .Q(acc_point_o[701]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][702] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][702]_srl3_n_0 ),
        .Q(acc_point_o[702]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][703] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][703]_srl3_n_0 ),
        .Q(acc_point_o[703]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][704] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][704]_srl3_n_0 ),
        .Q(acc_point_o[704]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][705] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][705]_srl3_n_0 ),
        .Q(acc_point_o[705]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][706] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][706]_srl3_n_0 ),
        .Q(acc_point_o[706]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][707] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][707]_srl3_n_0 ),
        .Q(acc_point_o[707]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][708] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][708]_srl3_n_0 ),
        .Q(acc_point_o[708]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][709] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][709]_srl3_n_0 ),
        .Q(acc_point_o[709]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][70] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][70]_srl3_n_0 ),
        .Q(acc_point_o[70]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][710] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][710]_srl3_n_0 ),
        .Q(acc_point_o[710]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][711] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][711]_srl3_n_0 ),
        .Q(acc_point_o[711]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][712] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][712]_srl3_n_0 ),
        .Q(acc_point_o[712]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][713] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][713]_srl3_n_0 ),
        .Q(acc_point_o[713]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][714] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][714]_srl3_n_0 ),
        .Q(acc_point_o[714]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][715] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][715]_srl3_n_0 ),
        .Q(acc_point_o[715]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][716] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][716]_srl3_n_0 ),
        .Q(acc_point_o[716]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][717] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][717]_srl3_n_0 ),
        .Q(acc_point_o[717]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][718] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][718]_srl3_n_0 ),
        .Q(acc_point_o[718]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][719] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][719]_srl3_n_0 ),
        .Q(acc_point_o[719]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][71] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][71]_srl3_n_0 ),
        .Q(acc_point_o[71]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][720] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][720]_srl3_n_0 ),
        .Q(acc_point_o[720]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][721] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][721]_srl3_n_0 ),
        .Q(acc_point_o[721]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][722] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][722]_srl3_n_0 ),
        .Q(acc_point_o[722]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][723] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][723]_srl3_n_0 ),
        .Q(acc_point_o[723]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][724] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][724]_srl3_n_0 ),
        .Q(acc_point_o[724]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][725] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][725]_srl3_n_0 ),
        .Q(acc_point_o[725]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][726] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][726]_srl3_n_0 ),
        .Q(acc_point_o[726]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][727] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][727]_srl3_n_0 ),
        .Q(acc_point_o[727]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][728] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][728]_srl3_n_0 ),
        .Q(acc_point_o[728]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][729] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][729]_srl3_n_0 ),
        .Q(acc_point_o[729]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][72] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][72]_srl3_n_0 ),
        .Q(acc_point_o[72]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][730] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][730]_srl3_n_0 ),
        .Q(acc_point_o[730]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][731] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][731]_srl3_n_0 ),
        .Q(acc_point_o[731]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][732] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][732]_srl3_n_0 ),
        .Q(acc_point_o[732]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][733] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][733]_srl3_n_0 ),
        .Q(acc_point_o[733]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][734] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][734]_srl3_n_0 ),
        .Q(acc_point_o[734]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][735] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][735]_srl3_n_0 ),
        .Q(acc_point_o[735]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][736] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][736]_srl3_n_0 ),
        .Q(acc_point_o[736]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][737] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][737]_srl3_n_0 ),
        .Q(acc_point_o[737]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][738] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][738]_srl3_n_0 ),
        .Q(acc_point_o[738]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][739] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][739]_srl3_n_0 ),
        .Q(acc_point_o[739]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][73] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][73]_srl3_n_0 ),
        .Q(acc_point_o[73]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][740] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][740]_srl3_n_0 ),
        .Q(acc_point_o[740]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][741] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][741]_srl3_n_0 ),
        .Q(acc_point_o[741]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][742] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][742]_srl3_n_0 ),
        .Q(acc_point_o[742]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][743] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][743]_srl3_n_0 ),
        .Q(acc_point_o[743]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][744] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][744]_srl3_n_0 ),
        .Q(acc_point_o[744]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][745] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][745]_srl3_n_0 ),
        .Q(acc_point_o[745]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][746] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][746]_srl3_n_0 ),
        .Q(acc_point_o[746]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][747] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][747]_srl3_n_0 ),
        .Q(acc_point_o[747]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][748] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][748]_srl3_n_0 ),
        .Q(acc_point_o[748]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][749] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][749]_srl3_n_0 ),
        .Q(acc_point_o[749]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][74] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][74]_srl3_n_0 ),
        .Q(acc_point_o[74]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][750] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][750]_srl3_n_0 ),
        .Q(acc_point_o[750]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][751] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][751]_srl3_n_0 ),
        .Q(acc_point_o[751]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][752] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][752]_srl3_n_0 ),
        .Q(acc_point_o[752]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][753] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][753]_srl3_n_0 ),
        .Q(acc_point_o[753]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][754] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][754]_srl3_n_0 ),
        .Q(acc_point_o[754]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][755] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][755]_srl3_n_0 ),
        .Q(acc_point_o[755]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][756] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][756]_srl3_n_0 ),
        .Q(acc_point_o[756]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][757] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][757]_srl3_n_0 ),
        .Q(acc_point_o[757]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][758] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][758]_srl3_n_0 ),
        .Q(acc_point_o[758]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][759] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][759]_srl3_n_0 ),
        .Q(acc_point_o[759]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][75] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][75]_srl3_n_0 ),
        .Q(acc_point_o[75]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][760] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][760]_srl3_n_0 ),
        .Q(acc_point_o[760]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][761] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][761]_srl3_n_0 ),
        .Q(acc_point_o[761]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][762] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][762]_srl3_n_0 ),
        .Q(acc_point_o[762]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][763] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][763]_srl3_n_0 ),
        .Q(acc_point_o[763]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][764] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][764]_srl3_n_0 ),
        .Q(acc_point_o[764]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][765] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][765]_srl3_n_0 ),
        .Q(acc_point_o[765]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][766] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][766]_srl3_n_0 ),
        .Q(acc_point_o[766]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][767] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][767]_srl3_n_0 ),
        .Q(acc_point_o[767]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][768] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][768]_srl3_n_0 ),
        .Q(acc_point_o[768]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][769] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][769]_srl3_n_0 ),
        .Q(acc_point_o[769]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][76] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][76]_srl3_n_0 ),
        .Q(acc_point_o[76]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][770] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][770]_srl3_n_0 ),
        .Q(acc_point_o[770]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][771] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][771]_srl3_n_0 ),
        .Q(acc_point_o[771]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][772] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][772]_srl3_n_0 ),
        .Q(acc_point_o[772]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][773] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][773]_srl3_n_0 ),
        .Q(acc_point_o[773]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][774] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][774]_srl3_n_0 ),
        .Q(acc_point_o[774]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][775] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][775]_srl3_n_0 ),
        .Q(acc_point_o[775]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][776] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][776]_srl3_n_0 ),
        .Q(acc_point_o[776]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][777] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][777]_srl3_n_0 ),
        .Q(acc_point_o[777]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][778] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][778]_srl3_n_0 ),
        .Q(acc_point_o[778]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][779] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][779]_srl3_n_0 ),
        .Q(acc_point_o[779]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][77] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][77]_srl3_n_0 ),
        .Q(acc_point_o[77]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][780] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][780]_srl3_n_0 ),
        .Q(acc_point_o[780]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][781] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][781]_srl3_n_0 ),
        .Q(acc_point_o[781]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][782] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][782]_srl3_n_0 ),
        .Q(acc_point_o[782]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][783] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][783]_srl3_n_0 ),
        .Q(acc_point_o[783]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][784] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][784]_srl3_n_0 ),
        .Q(acc_point_o[784]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][785] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][785]_srl3_n_0 ),
        .Q(acc_point_o[785]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][786] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][786]_srl3_n_0 ),
        .Q(acc_point_o[786]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][787] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][787]_srl3_n_0 ),
        .Q(acc_point_o[787]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][788] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][788]_srl3_n_0 ),
        .Q(acc_point_o[788]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][789] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][789]_srl3_n_0 ),
        .Q(acc_point_o[789]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][78] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][78]_srl3_n_0 ),
        .Q(acc_point_o[78]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][790] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][790]_srl3_n_0 ),
        .Q(acc_point_o[790]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][791] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][791]_srl3_n_0 ),
        .Q(acc_point_o[791]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][792] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][792]_srl3_n_0 ),
        .Q(acc_point_o[792]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][793] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][793]_srl3_n_0 ),
        .Q(acc_point_o[793]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][794] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][794]_srl3_n_0 ),
        .Q(acc_point_o[794]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][795] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][795]_srl3_n_0 ),
        .Q(acc_point_o[795]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][796] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][796]_srl3_n_0 ),
        .Q(acc_point_o[796]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][797] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][797]_srl3_n_0 ),
        .Q(acc_point_o[797]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][798] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][798]_srl3_n_0 ),
        .Q(acc_point_o[798]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][799] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][799]_srl3_n_0 ),
        .Q(acc_point_o[799]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][79] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][79]_srl3_n_0 ),
        .Q(acc_point_o[79]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][7]_srl3_n_0 ),
        .Q(acc_point_o[7]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][800] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][800]_srl3_n_0 ),
        .Q(acc_point_o[800]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][801] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][801]_srl3_n_0 ),
        .Q(acc_point_o[801]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][802] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][802]_srl3_n_0 ),
        .Q(acc_point_o[802]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][803] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][803]_srl3_n_0 ),
        .Q(acc_point_o[803]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][804] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][804]_srl3_n_0 ),
        .Q(acc_point_o[804]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][805] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][805]_srl3_n_0 ),
        .Q(acc_point_o[805]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][806] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][806]_srl3_n_0 ),
        .Q(acc_point_o[806]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][807] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][807]_srl3_n_0 ),
        .Q(acc_point_o[807]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][808] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][808]_srl3_n_0 ),
        .Q(acc_point_o[808]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][809] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][809]_srl3_n_0 ),
        .Q(acc_point_o[809]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][80] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][80]_srl3_n_0 ),
        .Q(acc_point_o[80]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][810] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][810]_srl3_n_0 ),
        .Q(acc_point_o[810]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][811] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][811]_srl3_n_0 ),
        .Q(acc_point_o[811]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][812] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][812]_srl3_n_0 ),
        .Q(acc_point_o[812]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][813] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][813]_srl3_n_0 ),
        .Q(acc_point_o[813]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][814] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][814]_srl3_n_0 ),
        .Q(acc_point_o[814]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][815] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][815]_srl3_n_0 ),
        .Q(acc_point_o[815]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][816] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][816]_srl3_n_0 ),
        .Q(acc_point_o[816]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][817] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][817]_srl3_n_0 ),
        .Q(acc_point_o[817]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][818] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][818]_srl3_n_0 ),
        .Q(acc_point_o[818]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][819] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][819]_srl3_n_0 ),
        .Q(acc_point_o[819]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][81] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][81]_srl3_n_0 ),
        .Q(acc_point_o[81]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][820] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][820]_srl3_n_0 ),
        .Q(acc_point_o[820]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][821] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][821]_srl3_n_0 ),
        .Q(acc_point_o[821]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][822] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][822]_srl3_n_0 ),
        .Q(acc_point_o[822]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][823] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][823]_srl3_n_0 ),
        .Q(acc_point_o[823]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][824] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][824]_srl3_n_0 ),
        .Q(acc_point_o[824]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][825] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][825]_srl3_n_0 ),
        .Q(acc_point_o[825]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][826] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][826]_srl3_n_0 ),
        .Q(acc_point_o[826]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][827] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][827]_srl3_n_0 ),
        .Q(acc_point_o[827]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][828] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][828]_srl3_n_0 ),
        .Q(acc_point_o[828]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][829] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][829]_srl3_n_0 ),
        .Q(acc_point_o[829]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][82] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][82]_srl3_n_0 ),
        .Q(acc_point_o[82]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][830] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][830]_srl3_n_0 ),
        .Q(acc_point_o[830]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][831] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][831]_srl3_n_0 ),
        .Q(acc_point_o[831]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][832] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][832]_srl3_n_0 ),
        .Q(acc_point_o[832]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][833] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][833]_srl3_n_0 ),
        .Q(acc_point_o[833]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][834] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][834]_srl3_n_0 ),
        .Q(acc_point_o[834]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][835] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][835]_srl3_n_0 ),
        .Q(acc_point_o[835]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][836] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][836]_srl3_n_0 ),
        .Q(acc_point_o[836]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][837] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][837]_srl3_n_0 ),
        .Q(acc_point_o[837]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][838] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][838]_srl3_n_0 ),
        .Q(acc_point_o[838]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][839] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][839]_srl3_n_0 ),
        .Q(acc_point_o[839]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][83] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][83]_srl3_n_0 ),
        .Q(acc_point_o[83]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][840] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][840]_srl3_n_0 ),
        .Q(acc_point_o[840]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][841] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][841]_srl3_n_0 ),
        .Q(acc_point_o[841]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][842] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][842]_srl3_n_0 ),
        .Q(acc_point_o[842]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][843] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][843]_srl3_n_0 ),
        .Q(acc_point_o[843]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][844] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][844]_srl3_n_0 ),
        .Q(acc_point_o[844]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][845] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][845]_srl3_n_0 ),
        .Q(acc_point_o[845]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][846] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][846]_srl3_n_0 ),
        .Q(acc_point_o[846]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][847] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][847]_srl3_n_0 ),
        .Q(acc_point_o[847]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][848] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][848]_srl3_n_0 ),
        .Q(acc_point_o[848]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][849] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][849]_srl3_n_0 ),
        .Q(acc_point_o[849]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][84] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][84]_srl3_n_0 ),
        .Q(acc_point_o[84]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][850] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][850]_srl3_n_0 ),
        .Q(acc_point_o[850]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][851] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][851]_srl3_n_0 ),
        .Q(acc_point_o[851]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][852] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][852]_srl3_n_0 ),
        .Q(acc_point_o[852]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][853] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][853]_srl3_n_0 ),
        .Q(acc_point_o[853]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][854] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][854]_srl3_n_0 ),
        .Q(acc_point_o[854]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][855] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][855]_srl3_n_0 ),
        .Q(acc_point_o[855]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][856] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][856]_srl3_n_0 ),
        .Q(acc_point_o[856]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][857] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][857]_srl3_n_0 ),
        .Q(acc_point_o[857]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][858] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][858]_srl3_n_0 ),
        .Q(acc_point_o[858]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][859] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][859]_srl3_n_0 ),
        .Q(acc_point_o[859]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][85] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][85]_srl3_n_0 ),
        .Q(acc_point_o[85]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][860] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][860]_srl3_n_0 ),
        .Q(acc_point_o[860]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][861] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][861]_srl3_n_0 ),
        .Q(acc_point_o[861]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][862] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][862]_srl3_n_0 ),
        .Q(acc_point_o[862]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][863] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][863]_srl3_n_0 ),
        .Q(acc_point_o[863]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][864] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][864]_srl3_n_0 ),
        .Q(acc_point_o[864]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][865] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][865]_srl3_n_0 ),
        .Q(acc_point_o[865]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][866] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][866]_srl3_n_0 ),
        .Q(acc_point_o[866]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][867] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][867]_srl3_n_0 ),
        .Q(acc_point_o[867]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][868] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][868]_srl3_n_0 ),
        .Q(acc_point_o[868]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][869] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][869]_srl3_n_0 ),
        .Q(acc_point_o[869]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][86] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][86]_srl3_n_0 ),
        .Q(acc_point_o[86]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][870] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][870]_srl3_n_0 ),
        .Q(acc_point_o[870]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][871] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][871]_srl3_n_0 ),
        .Q(acc_point_o[871]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][872] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][872]_srl3_n_0 ),
        .Q(acc_point_o[872]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][873] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][873]_srl3_n_0 ),
        .Q(acc_point_o[873]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][874] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][874]_srl3_n_0 ),
        .Q(acc_point_o[874]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][875] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][875]_srl3_n_0 ),
        .Q(acc_point_o[875]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][876] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][876]_srl3_n_0 ),
        .Q(acc_point_o[876]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][877] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][877]_srl3_n_0 ),
        .Q(acc_point_o[877]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][878] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][878]_srl3_n_0 ),
        .Q(acc_point_o[878]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][879] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][879]_srl3_n_0 ),
        .Q(acc_point_o[879]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][87] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][87]_srl3_n_0 ),
        .Q(acc_point_o[87]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][880] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][880]_srl3_n_0 ),
        .Q(acc_point_o[880]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][881] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][881]_srl3_n_0 ),
        .Q(acc_point_o[881]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][882] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][882]_srl3_n_0 ),
        .Q(acc_point_o[882]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][883] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][883]_srl3_n_0 ),
        .Q(acc_point_o[883]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][884] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][884]_srl3_n_0 ),
        .Q(acc_point_o[884]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][885] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][885]_srl3_n_0 ),
        .Q(acc_point_o[885]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][886] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][886]_srl3_n_0 ),
        .Q(acc_point_o[886]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][887] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][887]_srl3_n_0 ),
        .Q(acc_point_o[887]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][888] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][888]_srl3_n_0 ),
        .Q(acc_point_o[888]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][889] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][889]_srl3_n_0 ),
        .Q(acc_point_o[889]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][88] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][88]_srl3_n_0 ),
        .Q(acc_point_o[88]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][890] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][890]_srl3_n_0 ),
        .Q(acc_point_o[890]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][891] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][891]_srl3_n_0 ),
        .Q(acc_point_o[891]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][892] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][892]_srl3_n_0 ),
        .Q(acc_point_o[892]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][893] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][893]_srl3_n_0 ),
        .Q(acc_point_o[893]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][894] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][894]_srl3_n_0 ),
        .Q(acc_point_o[894]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][895] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][895]_srl3_n_0 ),
        .Q(acc_point_o[895]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][896] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][896]_srl3_n_0 ),
        .Q(acc_point_o[896]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][897] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][897]_srl3_n_0 ),
        .Q(acc_point_o[897]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][898] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][898]_srl3_n_0 ),
        .Q(acc_point_o[898]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][899] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][899]_srl3_n_0 ),
        .Q(acc_point_o[899]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][89] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][89]_srl3_n_0 ),
        .Q(acc_point_o[89]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][8]_srl3_n_0 ),
        .Q(acc_point_o[8]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][900] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][900]_srl3_n_0 ),
        .Q(acc_point_o[900]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][901] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][901]_srl3_n_0 ),
        .Q(acc_point_o[901]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][902] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][902]_srl3_n_0 ),
        .Q(acc_point_o[902]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][903] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][903]_srl3_n_0 ),
        .Q(acc_point_o[903]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][904] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][904]_srl3_n_0 ),
        .Q(acc_point_o[904]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][905] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][905]_srl3_n_0 ),
        .Q(acc_point_o[905]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][906] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][906]_srl3_n_0 ),
        .Q(acc_point_o[906]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][907] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][907]_srl3_n_0 ),
        .Q(acc_point_o[907]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][908] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][908]_srl3_n_0 ),
        .Q(acc_point_o[908]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][909] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][909]_srl3_n_0 ),
        .Q(acc_point_o[909]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][90] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][90]_srl3_n_0 ),
        .Q(acc_point_o[90]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][910] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][910]_srl3_n_0 ),
        .Q(acc_point_o[910]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][911] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][911]_srl3_n_0 ),
        .Q(acc_point_o[911]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][912] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][912]_srl3_n_0 ),
        .Q(acc_point_o[912]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][913] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][913]_srl3_n_0 ),
        .Q(acc_point_o[913]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][914] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][914]_srl3_n_0 ),
        .Q(acc_point_o[914]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][915] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][915]_srl3_n_0 ),
        .Q(acc_point_o[915]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][916] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][916]_srl3_n_0 ),
        .Q(acc_point_o[916]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][917] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][917]_srl3_n_0 ),
        .Q(acc_point_o[917]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][918] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][918]_srl3_n_0 ),
        .Q(acc_point_o[918]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][919] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][919]_srl3_n_0 ),
        .Q(acc_point_o[919]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][91] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][91]_srl3_n_0 ),
        .Q(acc_point_o[91]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][920] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][920]_srl3_n_0 ),
        .Q(acc_point_o[920]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][921] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][921]_srl3_n_0 ),
        .Q(acc_point_o[921]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][922] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][922]_srl3_n_0 ),
        .Q(acc_point_o[922]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][923] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][923]_srl3_n_0 ),
        .Q(acc_point_o[923]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][924] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][924]_srl3_n_0 ),
        .Q(acc_point_o[924]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][925] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][925]_srl3_n_0 ),
        .Q(acc_point_o[925]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][926] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][926]_srl3_n_0 ),
        .Q(acc_point_o[926]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][927] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][927]_srl3_n_0 ),
        .Q(acc_point_o[927]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][928] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][928]_srl3_n_0 ),
        .Q(acc_point_o[928]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][929] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][929]_srl3_n_0 ),
        .Q(acc_point_o[929]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][92] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][92]_srl3_n_0 ),
        .Q(acc_point_o[92]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][930] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][930]_srl3_n_0 ),
        .Q(acc_point_o[930]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][931] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][931]_srl3_n_0 ),
        .Q(acc_point_o[931]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][932] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][932]_srl3_n_0 ),
        .Q(acc_point_o[932]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][933] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][933]_srl3_n_0 ),
        .Q(acc_point_o[933]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][934] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][934]_srl3_n_0 ),
        .Q(acc_point_o[934]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][935] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][935]_srl3_n_0 ),
        .Q(acc_point_o[935]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][936] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][936]_srl3_n_0 ),
        .Q(acc_point_o[936]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][937] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][937]_srl3_n_0 ),
        .Q(acc_point_o[937]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][938] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][938]_srl3_n_0 ),
        .Q(acc_point_o[938]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][939] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][939]_srl3_n_0 ),
        .Q(acc_point_o[939]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][93] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][93]_srl3_n_0 ),
        .Q(acc_point_o[93]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][940] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][940]_srl3_n_0 ),
        .Q(acc_point_o[940]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][941] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][941]_srl3_n_0 ),
        .Q(acc_point_o[941]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][942] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][942]_srl3_n_0 ),
        .Q(acc_point_o[942]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][943] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][943]_srl3_n_0 ),
        .Q(acc_point_o[943]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][944] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][944]_srl3_n_0 ),
        .Q(acc_point_o[944]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][945] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][945]_srl3_n_0 ),
        .Q(acc_point_o[945]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][946] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][946]_srl3_n_0 ),
        .Q(acc_point_o[946]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][947] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][947]_srl3_n_0 ),
        .Q(acc_point_o[947]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][948] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][948]_srl3_n_0 ),
        .Q(acc_point_o[948]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][949] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][949]_srl3_n_0 ),
        .Q(acc_point_o[949]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][94] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][94]_srl3_n_0 ),
        .Q(acc_point_o[94]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][950] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][950]_srl3_n_0 ),
        .Q(acc_point_o[950]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][951] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][951]_srl3_n_0 ),
        .Q(acc_point_o[951]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][952] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][952]_srl3_n_0 ),
        .Q(acc_point_o[952]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][953] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][953]_srl3_n_0 ),
        .Q(acc_point_o[953]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][954] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][954]_srl3_n_0 ),
        .Q(acc_point_o[954]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][955] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][955]_srl3_n_0 ),
        .Q(acc_point_o[955]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][956] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][956]_srl3_n_0 ),
        .Q(acc_point_o[956]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][957] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][957]_srl3_n_0 ),
        .Q(acc_point_o[957]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][958] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][958]_srl3_n_0 ),
        .Q(acc_point_o[958]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][959] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][959]_srl3_n_0 ),
        .Q(acc_point_o[959]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][95] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][95]_srl3_n_0 ),
        .Q(acc_point_o[95]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][960] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][960]_srl3_n_0 ),
        .Q(acc_point_o[960]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][961] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][961]_srl3_n_0 ),
        .Q(acc_point_o[961]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][962] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][962]_srl3_n_0 ),
        .Q(acc_point_o[962]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][963] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][963]_srl3_n_0 ),
        .Q(acc_point_o[963]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][964] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][964]_srl3_n_0 ),
        .Q(acc_point_o[964]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][965] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][965]_srl3_n_0 ),
        .Q(acc_point_o[965]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][966] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][966]_srl3_n_0 ),
        .Q(acc_point_o[966]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][967] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][967]_srl3_n_0 ),
        .Q(acc_point_o[967]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][968] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][968]_srl3_n_0 ),
        .Q(acc_point_o[968]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][969] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][969]_srl3_n_0 ),
        .Q(acc_point_o[969]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][96] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][96]_srl3_n_0 ),
        .Q(acc_point_o[96]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][970] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][970]_srl3_n_0 ),
        .Q(acc_point_o[970]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][971] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][971]_srl3_n_0 ),
        .Q(acc_point_o[971]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][972] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][972]_srl3_n_0 ),
        .Q(acc_point_o[972]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][973] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][973]_srl3_n_0 ),
        .Q(acc_point_o[973]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][974] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][974]_srl3_n_0 ),
        .Q(acc_point_o[974]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][975] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][975]_srl3_n_0 ),
        .Q(acc_point_o[975]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][976] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][976]_srl3_n_0 ),
        .Q(acc_point_o[976]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][977] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][977]_srl3_n_0 ),
        .Q(acc_point_o[977]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][978] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][978]_srl3_n_0 ),
        .Q(acc_point_o[978]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][979] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][979]_srl3_n_0 ),
        .Q(acc_point_o[979]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][97] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][97]_srl3_n_0 ),
        .Q(acc_point_o[97]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][980] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][980]_srl3_n_0 ),
        .Q(acc_point_o[980]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][981] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][981]_srl3_n_0 ),
        .Q(acc_point_o[981]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][982] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][982]_srl3_n_0 ),
        .Q(acc_point_o[982]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][983] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][983]_srl3_n_0 ),
        .Q(acc_point_o[983]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][984] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][984]_srl3_n_0 ),
        .Q(acc_point_o[984]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][985] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][985]_srl3_n_0 ),
        .Q(acc_point_o[985]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][986] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][986]_srl3_n_0 ),
        .Q(acc_point_o[986]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][987] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][987]_srl3_n_0 ),
        .Q(acc_point_o[987]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][988] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][988]_srl3_n_0 ),
        .Q(acc_point_o[988]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][989] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][989]_srl3_n_0 ),
        .Q(acc_point_o[989]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][98] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][98]_srl3_n_0 ),
        .Q(acc_point_o[98]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][990] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][990]_srl3_n_0 ),
        .Q(acc_point_o[990]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][991] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][991]_srl3_n_0 ),
        .Q(acc_point_o[991]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][992] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][992]_srl3_n_0 ),
        .Q(acc_point_o[992]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][993] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][993]_srl3_n_0 ),
        .Q(acc_point_o[993]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][994] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][994]_srl3_n_0 ),
        .Q(acc_point_o[994]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][995] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][995]_srl3_n_0 ),
        .Q(acc_point_o[995]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][996] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][996]_srl3_n_0 ),
        .Q(acc_point_o[996]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][997] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][997]_srl3_n_0 ),
        .Q(acc_point_o[997]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][998] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][998]_srl3_n_0 ),
        .Q(acc_point_o[998]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][999] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][999]_srl3_n_0 ),
        .Q(acc_point_o[999]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][99] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][99]_srl3_n_0 ),
        .Q(acc_point_o[99]),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \DELAY_BLOCK[4].shift_array_reg[5][9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4][9]_srl3_n_0 ),
        .Q(acc_point_o[9]),
        .R(\<const0> ));
  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[0]),
        .Q(\shift_array_reg_n_0_[1][0] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1000] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1000]),
        .Q(\shift_array_reg_n_0_[1][1000] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1001] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1001]),
        .Q(\shift_array_reg_n_0_[1][1001] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1002] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1002]),
        .Q(\shift_array_reg_n_0_[1][1002] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1003] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1003]),
        .Q(\shift_array_reg_n_0_[1][1003] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1004] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1004]),
        .Q(\shift_array_reg_n_0_[1][1004] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1005] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1005]),
        .Q(\shift_array_reg_n_0_[1][1005] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1006] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1006]),
        .Q(\shift_array_reg_n_0_[1][1006] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1007] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1007]),
        .Q(\shift_array_reg_n_0_[1][1007] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1008] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1008]),
        .Q(\shift_array_reg_n_0_[1][1008] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1009] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1009]),
        .Q(\shift_array_reg_n_0_[1][1009] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][100] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[100]),
        .Q(\shift_array_reg_n_0_[1][100] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1010] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1010]),
        .Q(\shift_array_reg_n_0_[1][1010] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1011] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1011]),
        .Q(\shift_array_reg_n_0_[1][1011] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1012] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1012]),
        .Q(\shift_array_reg_n_0_[1][1012] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1013] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1013]),
        .Q(\shift_array_reg_n_0_[1][1013] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1014] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1014]),
        .Q(\shift_array_reg_n_0_[1][1014] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1015] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1015]),
        .Q(\shift_array_reg_n_0_[1][1015] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1016] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1016]),
        .Q(\shift_array_reg_n_0_[1][1016] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1017] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1017]),
        .Q(\shift_array_reg_n_0_[1][1017] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1018] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1018]),
        .Q(\shift_array_reg_n_0_[1][1018] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1019] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1019]),
        .Q(\shift_array_reg_n_0_[1][1019] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][101] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[101]),
        .Q(\shift_array_reg_n_0_[1][101] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1020] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1020]),
        .Q(\shift_array_reg_n_0_[1][1020] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1021] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1021]),
        .Q(\shift_array_reg_n_0_[1][1021] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1022] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1022]),
        .Q(\shift_array_reg_n_0_[1][1022] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1023] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1023]),
        .Q(\shift_array_reg_n_0_[1][1023] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1024] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1024]),
        .Q(\shift_array_reg_n_0_[1][1024] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1025] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1025]),
        .Q(\shift_array_reg_n_0_[1][1025] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1026] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1026]),
        .Q(\shift_array_reg_n_0_[1][1026] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1027] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1027]),
        .Q(\shift_array_reg_n_0_[1][1027] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1028] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1028]),
        .Q(\shift_array_reg_n_0_[1][1028] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1029] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1029]),
        .Q(\shift_array_reg_n_0_[1][1029] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][102] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[102]),
        .Q(\shift_array_reg_n_0_[1][102] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1030] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1030]),
        .Q(\shift_array_reg_n_0_[1][1030] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1031] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1031]),
        .Q(\shift_array_reg_n_0_[1][1031] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1032] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1032]),
        .Q(\shift_array_reg_n_0_[1][1032] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1033] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1033]),
        .Q(\shift_array_reg_n_0_[1][1033] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1034] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1034]),
        .Q(\shift_array_reg_n_0_[1][1034] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1035] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1035]),
        .Q(\shift_array_reg_n_0_[1][1035] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1036] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1036]),
        .Q(\shift_array_reg_n_0_[1][1036] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1037] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1037]),
        .Q(\shift_array_reg_n_0_[1][1037] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1038] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1038]),
        .Q(\shift_array_reg_n_0_[1][1038] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1039] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1039]),
        .Q(\shift_array_reg_n_0_[1][1039] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][103] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[103]),
        .Q(\shift_array_reg_n_0_[1][103] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1040] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1040]),
        .Q(\shift_array_reg_n_0_[1][1040] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1041] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1041]),
        .Q(\shift_array_reg_n_0_[1][1041] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1042] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1042]),
        .Q(\shift_array_reg_n_0_[1][1042] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1043] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1043]),
        .Q(\shift_array_reg_n_0_[1][1043] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1044] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1044]),
        .Q(\shift_array_reg_n_0_[1][1044] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1045] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1045]),
        .Q(\shift_array_reg_n_0_[1][1045] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1046] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1046]),
        .Q(\shift_array_reg_n_0_[1][1046] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1047] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1047]),
        .Q(\shift_array_reg_n_0_[1][1047] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1048] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1048]),
        .Q(\shift_array_reg_n_0_[1][1048] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1049] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1049]),
        .Q(\shift_array_reg_n_0_[1][1049] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][104] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[104]),
        .Q(\shift_array_reg_n_0_[1][104] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1050] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1050]),
        .Q(\shift_array_reg_n_0_[1][1050] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1051] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1051]),
        .Q(\shift_array_reg_n_0_[1][1051] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1052] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1052]),
        .Q(\shift_array_reg_n_0_[1][1052] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1053] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1053]),
        .Q(\shift_array_reg_n_0_[1][1053] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1054] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1054]),
        .Q(\shift_array_reg_n_0_[1][1054] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1055] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1055]),
        .Q(\shift_array_reg_n_0_[1][1055] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1056] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1056]),
        .Q(\shift_array_reg_n_0_[1][1056] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1057] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1057]),
        .Q(\shift_array_reg_n_0_[1][1057] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1058] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1058]),
        .Q(\shift_array_reg_n_0_[1][1058] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1059] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1059]),
        .Q(\shift_array_reg_n_0_[1][1059] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][105] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[105]),
        .Q(\shift_array_reg_n_0_[1][105] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1060] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1060]),
        .Q(\shift_array_reg_n_0_[1][1060] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1061] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1061]),
        .Q(\shift_array_reg_n_0_[1][1061] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1062] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1062]),
        .Q(\shift_array_reg_n_0_[1][1062] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1063] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1063]),
        .Q(\shift_array_reg_n_0_[1][1063] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1064] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1064]),
        .Q(\shift_array_reg_n_0_[1][1064] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1065] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1065]),
        .Q(\shift_array_reg_n_0_[1][1065] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1066] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1066]),
        .Q(\shift_array_reg_n_0_[1][1066] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1067] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1067]),
        .Q(\shift_array_reg_n_0_[1][1067] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1068] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1068]),
        .Q(\shift_array_reg_n_0_[1][1068] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1069] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1069]),
        .Q(\shift_array_reg_n_0_[1][1069] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][106] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[106]),
        .Q(\shift_array_reg_n_0_[1][106] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1070] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1070]),
        .Q(\shift_array_reg_n_0_[1][1070] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1071] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1071]),
        .Q(\shift_array_reg_n_0_[1][1071] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1072] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1072]),
        .Q(\shift_array_reg_n_0_[1][1072] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1073] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1073]),
        .Q(\shift_array_reg_n_0_[1][1073] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1074] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1074]),
        .Q(\shift_array_reg_n_0_[1][1074] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1075] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1075]),
        .Q(\shift_array_reg_n_0_[1][1075] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1076] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1076]),
        .Q(\shift_array_reg_n_0_[1][1076] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1077] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1077]),
        .Q(\shift_array_reg_n_0_[1][1077] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1078] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1078]),
        .Q(\shift_array_reg_n_0_[1][1078] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1079] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1079]),
        .Q(\shift_array_reg_n_0_[1][1079] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][107] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[107]),
        .Q(\shift_array_reg_n_0_[1][107] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1080] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1080]),
        .Q(\shift_array_reg_n_0_[1][1080] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1081] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1081]),
        .Q(\shift_array_reg_n_0_[1][1081] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1082] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1082]),
        .Q(\shift_array_reg_n_0_[1][1082] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1083] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1083]),
        .Q(\shift_array_reg_n_0_[1][1083] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1084] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1084]),
        .Q(\shift_array_reg_n_0_[1][1084] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1085] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1085]),
        .Q(\shift_array_reg_n_0_[1][1085] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1086] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1086]),
        .Q(\shift_array_reg_n_0_[1][1086] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1087] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1087]),
        .Q(\shift_array_reg_n_0_[1][1087] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1088] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1088]),
        .Q(\shift_array_reg_n_0_[1][1088] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1089] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1089]),
        .Q(\shift_array_reg_n_0_[1][1089] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][108] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[108]),
        .Q(\shift_array_reg_n_0_[1][108] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1090] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1090]),
        .Q(\shift_array_reg_n_0_[1][1090] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1091] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1091]),
        .Q(\shift_array_reg_n_0_[1][1091] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1092] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1092]),
        .Q(\shift_array_reg_n_0_[1][1092] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1093] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1093]),
        .Q(\shift_array_reg_n_0_[1][1093] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1094] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1094]),
        .Q(\shift_array_reg_n_0_[1][1094] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1095] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1095]),
        .Q(\shift_array_reg_n_0_[1][1095] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1096] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1096]),
        .Q(\shift_array_reg_n_0_[1][1096] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1097] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1097]),
        .Q(\shift_array_reg_n_0_[1][1097] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1098] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1098]),
        .Q(\shift_array_reg_n_0_[1][1098] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1099] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1099]),
        .Q(\shift_array_reg_n_0_[1][1099] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][109] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[109]),
        .Q(\shift_array_reg_n_0_[1][109] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[10]),
        .Q(\shift_array_reg_n_0_[1][10] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1100] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1100]),
        .Q(\shift_array_reg_n_0_[1][1100] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1101] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1101]),
        .Q(\shift_array_reg_n_0_[1][1101] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1102] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1102]),
        .Q(\shift_array_reg_n_0_[1][1102] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1103] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1103]),
        .Q(\shift_array_reg_n_0_[1][1103] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1104] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1104]),
        .Q(\shift_array_reg_n_0_[1][1104] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1105] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1105]),
        .Q(\shift_array_reg_n_0_[1][1105] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1106] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1106]),
        .Q(\shift_array_reg_n_0_[1][1106] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1107] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1107]),
        .Q(\shift_array_reg_n_0_[1][1107] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1108] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1108]),
        .Q(\shift_array_reg_n_0_[1][1108] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1109] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1109]),
        .Q(\shift_array_reg_n_0_[1][1109] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][110] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[110]),
        .Q(\shift_array_reg_n_0_[1][110] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1110] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1110]),
        .Q(\shift_array_reg_n_0_[1][1110] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1111] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1111]),
        .Q(\shift_array_reg_n_0_[1][1111] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1112] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1112]),
        .Q(\shift_array_reg_n_0_[1][1112] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1113] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1113]),
        .Q(\shift_array_reg_n_0_[1][1113] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1114] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1114]),
        .Q(\shift_array_reg_n_0_[1][1114] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1115] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1115]),
        .Q(\shift_array_reg_n_0_[1][1115] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1116] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1116]),
        .Q(\shift_array_reg_n_0_[1][1116] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1117] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1117]),
        .Q(\shift_array_reg_n_0_[1][1117] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1118] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1118]),
        .Q(\shift_array_reg_n_0_[1][1118] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1119] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1119]),
        .Q(\shift_array_reg_n_0_[1][1119] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][111] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[111]),
        .Q(\shift_array_reg_n_0_[1][111] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1120] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1120]),
        .Q(\shift_array_reg_n_0_[1][1120] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1121] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1121]),
        .Q(\shift_array_reg_n_0_[1][1121] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1122] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1122]),
        .Q(\shift_array_reg_n_0_[1][1122] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1123] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1123]),
        .Q(\shift_array_reg_n_0_[1][1123] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1124] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1124]),
        .Q(\shift_array_reg_n_0_[1][1124] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1125] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1125]),
        .Q(\shift_array_reg_n_0_[1][1125] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1126] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1126]),
        .Q(\shift_array_reg_n_0_[1][1126] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1127] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1127]),
        .Q(\shift_array_reg_n_0_[1][1127] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1128] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1128]),
        .Q(\shift_array_reg_n_0_[1][1128] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1129] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1129]),
        .Q(\shift_array_reg_n_0_[1][1129] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][112] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[112]),
        .Q(\shift_array_reg_n_0_[1][112] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1130] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1130]),
        .Q(\shift_array_reg_n_0_[1][1130] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1131] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1131]),
        .Q(\shift_array_reg_n_0_[1][1131] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1132] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1132]),
        .Q(\shift_array_reg_n_0_[1][1132] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1133] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1133]),
        .Q(\shift_array_reg_n_0_[1][1133] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1134] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1134]),
        .Q(\shift_array_reg_n_0_[1][1134] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1135] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1135]),
        .Q(\shift_array_reg_n_0_[1][1135] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1136] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1136]),
        .Q(\shift_array_reg_n_0_[1][1136] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1137] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1137]),
        .Q(\shift_array_reg_n_0_[1][1137] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1138] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1138]),
        .Q(\shift_array_reg_n_0_[1][1138] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1139] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1139]),
        .Q(\shift_array_reg_n_0_[1][1139] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][113] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[113]),
        .Q(\shift_array_reg_n_0_[1][113] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1140] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1140]),
        .Q(\shift_array_reg_n_0_[1][1140] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1141] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1141]),
        .Q(\shift_array_reg_n_0_[1][1141] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1142] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1142]),
        .Q(\shift_array_reg_n_0_[1][1142] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1143] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1143]),
        .Q(\shift_array_reg_n_0_[1][1143] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1144] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1144]),
        .Q(\shift_array_reg_n_0_[1][1144] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1145] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1145]),
        .Q(\shift_array_reg_n_0_[1][1145] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1146] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1146]),
        .Q(\shift_array_reg_n_0_[1][1146] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1147] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1147]),
        .Q(\shift_array_reg_n_0_[1][1147] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1148] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1148]),
        .Q(\shift_array_reg_n_0_[1][1148] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1149] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1149]),
        .Q(\shift_array_reg_n_0_[1][1149] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][114] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[114]),
        .Q(\shift_array_reg_n_0_[1][114] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1150] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1150]),
        .Q(\shift_array_reg_n_0_[1][1150] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1151] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1151]),
        .Q(\shift_array_reg_n_0_[1][1151] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1152] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1152]),
        .Q(\shift_array_reg_n_0_[1][1152] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1153] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1153]),
        .Q(\shift_array_reg_n_0_[1][1153] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1154] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1154]),
        .Q(\shift_array_reg_n_0_[1][1154] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1155] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1155]),
        .Q(\shift_array_reg_n_0_[1][1155] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1156] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1156]),
        .Q(\shift_array_reg_n_0_[1][1156] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1157] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1157]),
        .Q(\shift_array_reg_n_0_[1][1157] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1158] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1158]),
        .Q(\shift_array_reg_n_0_[1][1158] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1159] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1159]),
        .Q(\shift_array_reg_n_0_[1][1159] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][115] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[115]),
        .Q(\shift_array_reg_n_0_[1][115] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1160] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1160]),
        .Q(\shift_array_reg_n_0_[1][1160] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1161] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1161]),
        .Q(\shift_array_reg_n_0_[1][1161] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1162] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1162]),
        .Q(\shift_array_reg_n_0_[1][1162] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1163] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1163]),
        .Q(\shift_array_reg_n_0_[1][1163] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][116] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[116]),
        .Q(\shift_array_reg_n_0_[1][116] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][117] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[117]),
        .Q(\shift_array_reg_n_0_[1][117] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][118] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[118]),
        .Q(\shift_array_reg_n_0_[1][118] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][119] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[119]),
        .Q(\shift_array_reg_n_0_[1][119] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[11]),
        .Q(\shift_array_reg_n_0_[1][11] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][120] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[120]),
        .Q(\shift_array_reg_n_0_[1][120] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][121] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[121]),
        .Q(\shift_array_reg_n_0_[1][121] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][122] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[122]),
        .Q(\shift_array_reg_n_0_[1][122] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][123] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[123]),
        .Q(\shift_array_reg_n_0_[1][123] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][124] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[124]),
        .Q(\shift_array_reg_n_0_[1][124] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][125] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[125]),
        .Q(\shift_array_reg_n_0_[1][125] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][126] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[126]),
        .Q(\shift_array_reg_n_0_[1][126] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][127] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[127]),
        .Q(\shift_array_reg_n_0_[1][127] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][128] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[128]),
        .Q(\shift_array_reg_n_0_[1][128] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][129] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[129]),
        .Q(\shift_array_reg_n_0_[1][129] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[12]),
        .Q(\shift_array_reg_n_0_[1][12] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][130] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[130]),
        .Q(\shift_array_reg_n_0_[1][130] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][131] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[131]),
        .Q(\shift_array_reg_n_0_[1][131] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][132] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[132]),
        .Q(\shift_array_reg_n_0_[1][132] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][133] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[133]),
        .Q(\shift_array_reg_n_0_[1][133] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][134] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[134]),
        .Q(\shift_array_reg_n_0_[1][134] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][135] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[135]),
        .Q(\shift_array_reg_n_0_[1][135] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][136] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[136]),
        .Q(\shift_array_reg_n_0_[1][136] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][137] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[137]),
        .Q(\shift_array_reg_n_0_[1][137] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][138] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[138]),
        .Q(\shift_array_reg_n_0_[1][138] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][139] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[139]),
        .Q(\shift_array_reg_n_0_[1][139] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[13]),
        .Q(\shift_array_reg_n_0_[1][13] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][140] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[140]),
        .Q(\shift_array_reg_n_0_[1][140] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][141] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[141]),
        .Q(\shift_array_reg_n_0_[1][141] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][142] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[142]),
        .Q(\shift_array_reg_n_0_[1][142] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][143] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[143]),
        .Q(\shift_array_reg_n_0_[1][143] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][144] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[144]),
        .Q(\shift_array_reg_n_0_[1][144] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][145] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[145]),
        .Q(\shift_array_reg_n_0_[1][145] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][146] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[146]),
        .Q(\shift_array_reg_n_0_[1][146] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][147] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[147]),
        .Q(\shift_array_reg_n_0_[1][147] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][148] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[148]),
        .Q(\shift_array_reg_n_0_[1][148] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][149] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[149]),
        .Q(\shift_array_reg_n_0_[1][149] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[14]),
        .Q(\shift_array_reg_n_0_[1][14] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][150] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[150]),
        .Q(\shift_array_reg_n_0_[1][150] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][151] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[151]),
        .Q(\shift_array_reg_n_0_[1][151] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][152] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[152]),
        .Q(\shift_array_reg_n_0_[1][152] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][153] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[153]),
        .Q(\shift_array_reg_n_0_[1][153] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][154] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[154]),
        .Q(\shift_array_reg_n_0_[1][154] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][155] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[155]),
        .Q(\shift_array_reg_n_0_[1][155] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][156] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[156]),
        .Q(\shift_array_reg_n_0_[1][156] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][157] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[157]),
        .Q(\shift_array_reg_n_0_[1][157] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][158] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[158]),
        .Q(\shift_array_reg_n_0_[1][158] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][159] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[159]),
        .Q(\shift_array_reg_n_0_[1][159] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[15]),
        .Q(\shift_array_reg_n_0_[1][15] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][160] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[160]),
        .Q(\shift_array_reg_n_0_[1][160] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][161] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[161]),
        .Q(\shift_array_reg_n_0_[1][161] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][162] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[162]),
        .Q(\shift_array_reg_n_0_[1][162] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][163] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[163]),
        .Q(\shift_array_reg_n_0_[1][163] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][164] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[164]),
        .Q(\shift_array_reg_n_0_[1][164] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][165] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[165]),
        .Q(\shift_array_reg_n_0_[1][165] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][166] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[166]),
        .Q(\shift_array_reg_n_0_[1][166] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][167] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[167]),
        .Q(\shift_array_reg_n_0_[1][167] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][168] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[168]),
        .Q(\shift_array_reg_n_0_[1][168] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][169] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[169]),
        .Q(\shift_array_reg_n_0_[1][169] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[16]),
        .Q(\shift_array_reg_n_0_[1][16] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][170] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[170]),
        .Q(\shift_array_reg_n_0_[1][170] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][171] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[171]),
        .Q(\shift_array_reg_n_0_[1][171] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][172] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[172]),
        .Q(\shift_array_reg_n_0_[1][172] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][173] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[173]),
        .Q(\shift_array_reg_n_0_[1][173] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][174] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[174]),
        .Q(\shift_array_reg_n_0_[1][174] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][175] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[175]),
        .Q(\shift_array_reg_n_0_[1][175] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][176] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[176]),
        .Q(\shift_array_reg_n_0_[1][176] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][177] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[177]),
        .Q(\shift_array_reg_n_0_[1][177] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][178] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[178]),
        .Q(\shift_array_reg_n_0_[1][178] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][179] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[179]),
        .Q(\shift_array_reg_n_0_[1][179] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[17]),
        .Q(\shift_array_reg_n_0_[1][17] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][180] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[180]),
        .Q(\shift_array_reg_n_0_[1][180] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][181] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[181]),
        .Q(\shift_array_reg_n_0_[1][181] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][182] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[182]),
        .Q(\shift_array_reg_n_0_[1][182] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][183] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[183]),
        .Q(\shift_array_reg_n_0_[1][183] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][184] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[184]),
        .Q(\shift_array_reg_n_0_[1][184] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][185] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[185]),
        .Q(\shift_array_reg_n_0_[1][185] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][186] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[186]),
        .Q(\shift_array_reg_n_0_[1][186] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][187] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[187]),
        .Q(\shift_array_reg_n_0_[1][187] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][188] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[188]),
        .Q(\shift_array_reg_n_0_[1][188] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][189] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[189]),
        .Q(\shift_array_reg_n_0_[1][189] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[18]),
        .Q(\shift_array_reg_n_0_[1][18] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][190] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[190]),
        .Q(\shift_array_reg_n_0_[1][190] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][191] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[191]),
        .Q(\shift_array_reg_n_0_[1][191] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][192] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[192]),
        .Q(\shift_array_reg_n_0_[1][192] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][193] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[193]),
        .Q(\shift_array_reg_n_0_[1][193] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][194] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[194]),
        .Q(\shift_array_reg_n_0_[1][194] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][195] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[195]),
        .Q(\shift_array_reg_n_0_[1][195] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][196] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[196]),
        .Q(\shift_array_reg_n_0_[1][196] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][197] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[197]),
        .Q(\shift_array_reg_n_0_[1][197] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][198] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[198]),
        .Q(\shift_array_reg_n_0_[1][198] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][199] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[199]),
        .Q(\shift_array_reg_n_0_[1][199] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[19]),
        .Q(\shift_array_reg_n_0_[1][19] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[1]),
        .Q(\shift_array_reg_n_0_[1][1] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][200] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[200]),
        .Q(\shift_array_reg_n_0_[1][200] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][201] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[201]),
        .Q(\shift_array_reg_n_0_[1][201] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][202] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[202]),
        .Q(\shift_array_reg_n_0_[1][202] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][203] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[203]),
        .Q(\shift_array_reg_n_0_[1][203] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][204] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[204]),
        .Q(\shift_array_reg_n_0_[1][204] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][205] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[205]),
        .Q(\shift_array_reg_n_0_[1][205] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][206] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[206]),
        .Q(\shift_array_reg_n_0_[1][206] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][207] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[207]),
        .Q(\shift_array_reg_n_0_[1][207] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][208] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[208]),
        .Q(\shift_array_reg_n_0_[1][208] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][209] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[209]),
        .Q(\shift_array_reg_n_0_[1][209] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[20]),
        .Q(\shift_array_reg_n_0_[1][20] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][210] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[210]),
        .Q(\shift_array_reg_n_0_[1][210] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][211] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[211]),
        .Q(\shift_array_reg_n_0_[1][211] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][212] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[212]),
        .Q(\shift_array_reg_n_0_[1][212] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][213] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[213]),
        .Q(\shift_array_reg_n_0_[1][213] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][214] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[214]),
        .Q(\shift_array_reg_n_0_[1][214] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][215] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[215]),
        .Q(\shift_array_reg_n_0_[1][215] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][216] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[216]),
        .Q(\shift_array_reg_n_0_[1][216] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][217] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[217]),
        .Q(\shift_array_reg_n_0_[1][217] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][218] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[218]),
        .Q(\shift_array_reg_n_0_[1][218] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][219] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[219]),
        .Q(\shift_array_reg_n_0_[1][219] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[21]),
        .Q(\shift_array_reg_n_0_[1][21] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][220] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[220]),
        .Q(\shift_array_reg_n_0_[1][220] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][221] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[221]),
        .Q(\shift_array_reg_n_0_[1][221] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][222] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[222]),
        .Q(\shift_array_reg_n_0_[1][222] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][223] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[223]),
        .Q(\shift_array_reg_n_0_[1][223] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][224] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[224]),
        .Q(\shift_array_reg_n_0_[1][224] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][225] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[225]),
        .Q(\shift_array_reg_n_0_[1][225] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][226] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[226]),
        .Q(\shift_array_reg_n_0_[1][226] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][227] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[227]),
        .Q(\shift_array_reg_n_0_[1][227] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][228] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[228]),
        .Q(\shift_array_reg_n_0_[1][228] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][229] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[229]),
        .Q(\shift_array_reg_n_0_[1][229] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[22]),
        .Q(\shift_array_reg_n_0_[1][22] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][230] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[230]),
        .Q(\shift_array_reg_n_0_[1][230] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][231] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[231]),
        .Q(\shift_array_reg_n_0_[1][231] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][232] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[232]),
        .Q(\shift_array_reg_n_0_[1][232] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][233] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[233]),
        .Q(\shift_array_reg_n_0_[1][233] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][234] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[234]),
        .Q(\shift_array_reg_n_0_[1][234] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][235] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[235]),
        .Q(\shift_array_reg_n_0_[1][235] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][236] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[236]),
        .Q(\shift_array_reg_n_0_[1][236] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][237] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[237]),
        .Q(\shift_array_reg_n_0_[1][237] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][238] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[238]),
        .Q(\shift_array_reg_n_0_[1][238] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][239] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[239]),
        .Q(\shift_array_reg_n_0_[1][239] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[23]),
        .Q(\shift_array_reg_n_0_[1][23] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][240] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[240]),
        .Q(\shift_array_reg_n_0_[1][240] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][241] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[241]),
        .Q(\shift_array_reg_n_0_[1][241] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][242] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[242]),
        .Q(\shift_array_reg_n_0_[1][242] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][243] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[243]),
        .Q(\shift_array_reg_n_0_[1][243] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][244] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[244]),
        .Q(\shift_array_reg_n_0_[1][244] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][245] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[245]),
        .Q(\shift_array_reg_n_0_[1][245] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][246] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[246]),
        .Q(\shift_array_reg_n_0_[1][246] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][247] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[247]),
        .Q(\shift_array_reg_n_0_[1][247] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][248] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[248]),
        .Q(\shift_array_reg_n_0_[1][248] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][249] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[249]),
        .Q(\shift_array_reg_n_0_[1][249] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[24]),
        .Q(\shift_array_reg_n_0_[1][24] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][250] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[250]),
        .Q(\shift_array_reg_n_0_[1][250] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][251] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[251]),
        .Q(\shift_array_reg_n_0_[1][251] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][252] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[252]),
        .Q(\shift_array_reg_n_0_[1][252] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][253] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[253]),
        .Q(\shift_array_reg_n_0_[1][253] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][254] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[254]),
        .Q(\shift_array_reg_n_0_[1][254] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][255] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[255]),
        .Q(\shift_array_reg_n_0_[1][255] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][256] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[256]),
        .Q(\shift_array_reg_n_0_[1][256] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][257] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[257]),
        .Q(\shift_array_reg_n_0_[1][257] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][258] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[258]),
        .Q(\shift_array_reg_n_0_[1][258] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][259] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[259]),
        .Q(\shift_array_reg_n_0_[1][259] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[25]),
        .Q(\shift_array_reg_n_0_[1][25] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][260] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[260]),
        .Q(\shift_array_reg_n_0_[1][260] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][261] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[261]),
        .Q(\shift_array_reg_n_0_[1][261] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][262] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[262]),
        .Q(\shift_array_reg_n_0_[1][262] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][263] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[263]),
        .Q(\shift_array_reg_n_0_[1][263] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][264] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[264]),
        .Q(\shift_array_reg_n_0_[1][264] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][265] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[265]),
        .Q(\shift_array_reg_n_0_[1][265] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][266] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[266]),
        .Q(\shift_array_reg_n_0_[1][266] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][267] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[267]),
        .Q(\shift_array_reg_n_0_[1][267] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][268] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[268]),
        .Q(\shift_array_reg_n_0_[1][268] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][269] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[269]),
        .Q(\shift_array_reg_n_0_[1][269] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[26]),
        .Q(\shift_array_reg_n_0_[1][26] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][270] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[270]),
        .Q(\shift_array_reg_n_0_[1][270] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][271] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[271]),
        .Q(\shift_array_reg_n_0_[1][271] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][272] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[272]),
        .Q(\shift_array_reg_n_0_[1][272] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][273] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[273]),
        .Q(\shift_array_reg_n_0_[1][273] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][274] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[274]),
        .Q(\shift_array_reg_n_0_[1][274] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][275] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[275]),
        .Q(\shift_array_reg_n_0_[1][275] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][276] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[276]),
        .Q(\shift_array_reg_n_0_[1][276] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][277] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[277]),
        .Q(\shift_array_reg_n_0_[1][277] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][278] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[278]),
        .Q(\shift_array_reg_n_0_[1][278] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][279] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[279]),
        .Q(\shift_array_reg_n_0_[1][279] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[27]),
        .Q(\shift_array_reg_n_0_[1][27] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][280] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[280]),
        .Q(\shift_array_reg_n_0_[1][280] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][281] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[281]),
        .Q(\shift_array_reg_n_0_[1][281] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][282] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[282]),
        .Q(\shift_array_reg_n_0_[1][282] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][283] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[283]),
        .Q(\shift_array_reg_n_0_[1][283] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][284] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[284]),
        .Q(\shift_array_reg_n_0_[1][284] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][285] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[285]),
        .Q(\shift_array_reg_n_0_[1][285] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][286] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[286]),
        .Q(\shift_array_reg_n_0_[1][286] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][287] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[287]),
        .Q(\shift_array_reg_n_0_[1][287] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][288] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[288]),
        .Q(\shift_array_reg_n_0_[1][288] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][289] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[289]),
        .Q(\shift_array_reg_n_0_[1][289] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[28]),
        .Q(\shift_array_reg_n_0_[1][28] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][290] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[290]),
        .Q(\shift_array_reg_n_0_[1][290] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][291] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[291]),
        .Q(\shift_array_reg_n_0_[1][291] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][292] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[292]),
        .Q(\shift_array_reg_n_0_[1][292] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][293] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[293]),
        .Q(\shift_array_reg_n_0_[1][293] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][294] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[294]),
        .Q(\shift_array_reg_n_0_[1][294] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][295] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[295]),
        .Q(\shift_array_reg_n_0_[1][295] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][296] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[296]),
        .Q(\shift_array_reg_n_0_[1][296] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][297] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[297]),
        .Q(\shift_array_reg_n_0_[1][297] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][298] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[298]),
        .Q(\shift_array_reg_n_0_[1][298] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][299] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[299]),
        .Q(\shift_array_reg_n_0_[1][299] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[29]),
        .Q(\shift_array_reg_n_0_[1][29] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[2]),
        .Q(\shift_array_reg_n_0_[1][2] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][300] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[300]),
        .Q(\shift_array_reg_n_0_[1][300] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][301] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[301]),
        .Q(\shift_array_reg_n_0_[1][301] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][302] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[302]),
        .Q(\shift_array_reg_n_0_[1][302] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][303] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[303]),
        .Q(\shift_array_reg_n_0_[1][303] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][304] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[304]),
        .Q(\shift_array_reg_n_0_[1][304] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][305] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[305]),
        .Q(\shift_array_reg_n_0_[1][305] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][306] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[306]),
        .Q(\shift_array_reg_n_0_[1][306] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][307] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[307]),
        .Q(\shift_array_reg_n_0_[1][307] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][308] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[308]),
        .Q(\shift_array_reg_n_0_[1][308] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][309] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[309]),
        .Q(\shift_array_reg_n_0_[1][309] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[30]),
        .Q(\shift_array_reg_n_0_[1][30] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][310] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[310]),
        .Q(\shift_array_reg_n_0_[1][310] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][311] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[311]),
        .Q(\shift_array_reg_n_0_[1][311] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][312] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[312]),
        .Q(\shift_array_reg_n_0_[1][312] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][313] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[313]),
        .Q(\shift_array_reg_n_0_[1][313] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][314] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[314]),
        .Q(\shift_array_reg_n_0_[1][314] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][315] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[315]),
        .Q(\shift_array_reg_n_0_[1][315] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][316] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[316]),
        .Q(\shift_array_reg_n_0_[1][316] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][317] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[317]),
        .Q(\shift_array_reg_n_0_[1][317] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][318] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[318]),
        .Q(\shift_array_reg_n_0_[1][318] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][319] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[319]),
        .Q(\shift_array_reg_n_0_[1][319] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[31]),
        .Q(\shift_array_reg_n_0_[1][31] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][320] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[320]),
        .Q(\shift_array_reg_n_0_[1][320] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][321] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[321]),
        .Q(\shift_array_reg_n_0_[1][321] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][322] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[322]),
        .Q(\shift_array_reg_n_0_[1][322] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][323] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[323]),
        .Q(\shift_array_reg_n_0_[1][323] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][324] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[324]),
        .Q(\shift_array_reg_n_0_[1][324] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][325] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[325]),
        .Q(\shift_array_reg_n_0_[1][325] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][326] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[326]),
        .Q(\shift_array_reg_n_0_[1][326] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][327] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[327]),
        .Q(\shift_array_reg_n_0_[1][327] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][328] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[328]),
        .Q(\shift_array_reg_n_0_[1][328] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][329] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[329]),
        .Q(\shift_array_reg_n_0_[1][329] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][32] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[32]),
        .Q(\shift_array_reg_n_0_[1][32] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][330] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[330]),
        .Q(\shift_array_reg_n_0_[1][330] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][331] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[331]),
        .Q(\shift_array_reg_n_0_[1][331] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][332] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[332]),
        .Q(\shift_array_reg_n_0_[1][332] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][333] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[333]),
        .Q(\shift_array_reg_n_0_[1][333] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][334] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[334]),
        .Q(\shift_array_reg_n_0_[1][334] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][335] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[335]),
        .Q(\shift_array_reg_n_0_[1][335] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][336] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[336]),
        .Q(\shift_array_reg_n_0_[1][336] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][337] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[337]),
        .Q(\shift_array_reg_n_0_[1][337] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][338] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[338]),
        .Q(\shift_array_reg_n_0_[1][338] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][339] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[339]),
        .Q(\shift_array_reg_n_0_[1][339] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][33] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[33]),
        .Q(\shift_array_reg_n_0_[1][33] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][340] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[340]),
        .Q(\shift_array_reg_n_0_[1][340] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][341] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[341]),
        .Q(\shift_array_reg_n_0_[1][341] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][342] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[342]),
        .Q(\shift_array_reg_n_0_[1][342] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][343] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[343]),
        .Q(\shift_array_reg_n_0_[1][343] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][344] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[344]),
        .Q(\shift_array_reg_n_0_[1][344] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][345] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[345]),
        .Q(\shift_array_reg_n_0_[1][345] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][346] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[346]),
        .Q(\shift_array_reg_n_0_[1][346] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][347] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[347]),
        .Q(\shift_array_reg_n_0_[1][347] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][348] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[348]),
        .Q(\shift_array_reg_n_0_[1][348] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][349] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[349]),
        .Q(\shift_array_reg_n_0_[1][349] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][34] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[34]),
        .Q(\shift_array_reg_n_0_[1][34] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][350] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[350]),
        .Q(\shift_array_reg_n_0_[1][350] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][351] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[351]),
        .Q(\shift_array_reg_n_0_[1][351] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][352] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[352]),
        .Q(\shift_array_reg_n_0_[1][352] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][353] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[353]),
        .Q(\shift_array_reg_n_0_[1][353] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][354] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[354]),
        .Q(\shift_array_reg_n_0_[1][354] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][355] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[355]),
        .Q(\shift_array_reg_n_0_[1][355] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][356] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[356]),
        .Q(\shift_array_reg_n_0_[1][356] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][357] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[357]),
        .Q(\shift_array_reg_n_0_[1][357] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][358] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[358]),
        .Q(\shift_array_reg_n_0_[1][358] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][359] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[359]),
        .Q(\shift_array_reg_n_0_[1][359] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][35] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[35]),
        .Q(\shift_array_reg_n_0_[1][35] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][360] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[360]),
        .Q(\shift_array_reg_n_0_[1][360] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][361] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[361]),
        .Q(\shift_array_reg_n_0_[1][361] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][362] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[362]),
        .Q(\shift_array_reg_n_0_[1][362] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][363] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[363]),
        .Q(\shift_array_reg_n_0_[1][363] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][364] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[364]),
        .Q(\shift_array_reg_n_0_[1][364] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][365] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[365]),
        .Q(\shift_array_reg_n_0_[1][365] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][366] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[366]),
        .Q(\shift_array_reg_n_0_[1][366] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][367] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[367]),
        .Q(\shift_array_reg_n_0_[1][367] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][368] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[368]),
        .Q(\shift_array_reg_n_0_[1][368] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][369] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[369]),
        .Q(\shift_array_reg_n_0_[1][369] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][36] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[36]),
        .Q(\shift_array_reg_n_0_[1][36] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][370] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[370]),
        .Q(\shift_array_reg_n_0_[1][370] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][371] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[371]),
        .Q(\shift_array_reg_n_0_[1][371] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][372] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[372]),
        .Q(\shift_array_reg_n_0_[1][372] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][373] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[373]),
        .Q(\shift_array_reg_n_0_[1][373] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][374] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[374]),
        .Q(\shift_array_reg_n_0_[1][374] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][375] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[375]),
        .Q(\shift_array_reg_n_0_[1][375] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][376] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[376]),
        .Q(\shift_array_reg_n_0_[1][376] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][377] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[377]),
        .Q(\shift_array_reg_n_0_[1][377] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][378] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[378]),
        .Q(\shift_array_reg_n_0_[1][378] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][379] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[379]),
        .Q(\shift_array_reg_n_0_[1][379] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][37] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[37]),
        .Q(\shift_array_reg_n_0_[1][37] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][380] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[380]),
        .Q(\shift_array_reg_n_0_[1][380] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][381] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[381]),
        .Q(\shift_array_reg_n_0_[1][381] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][382] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[382]),
        .Q(\shift_array_reg_n_0_[1][382] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][383] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[383]),
        .Q(\shift_array_reg_n_0_[1][383] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][384] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[384]),
        .Q(\shift_array_reg_n_0_[1][384] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][385] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[385]),
        .Q(\shift_array_reg_n_0_[1][385] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][386] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[386]),
        .Q(\shift_array_reg_n_0_[1][386] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][387] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[387]),
        .Q(\shift_array_reg_n_0_[1][387] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][388] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[388]),
        .Q(\shift_array_reg_n_0_[1][388] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][389] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[389]),
        .Q(\shift_array_reg_n_0_[1][389] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][38] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[38]),
        .Q(\shift_array_reg_n_0_[1][38] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][390] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[390]),
        .Q(\shift_array_reg_n_0_[1][390] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][391] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[391]),
        .Q(\shift_array_reg_n_0_[1][391] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][392] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[392]),
        .Q(\shift_array_reg_n_0_[1][392] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][393] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[393]),
        .Q(\shift_array_reg_n_0_[1][393] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][394] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[394]),
        .Q(\shift_array_reg_n_0_[1][394] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][395] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[395]),
        .Q(\shift_array_reg_n_0_[1][395] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][396] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[396]),
        .Q(\shift_array_reg_n_0_[1][396] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][397] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[397]),
        .Q(\shift_array_reg_n_0_[1][397] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][398] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[398]),
        .Q(\shift_array_reg_n_0_[1][398] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][399] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[399]),
        .Q(\shift_array_reg_n_0_[1][399] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][39] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[39]),
        .Q(\shift_array_reg_n_0_[1][39] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[3]),
        .Q(\shift_array_reg_n_0_[1][3] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][400] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[400]),
        .Q(\shift_array_reg_n_0_[1][400] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][401] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[401]),
        .Q(\shift_array_reg_n_0_[1][401] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][402] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[402]),
        .Q(\shift_array_reg_n_0_[1][402] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][403] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[403]),
        .Q(\shift_array_reg_n_0_[1][403] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][404] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[404]),
        .Q(\shift_array_reg_n_0_[1][404] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][405] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[405]),
        .Q(\shift_array_reg_n_0_[1][405] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][406] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[406]),
        .Q(\shift_array_reg_n_0_[1][406] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][407] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[407]),
        .Q(\shift_array_reg_n_0_[1][407] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][408] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[408]),
        .Q(\shift_array_reg_n_0_[1][408] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][409] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[409]),
        .Q(\shift_array_reg_n_0_[1][409] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][40] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[40]),
        .Q(\shift_array_reg_n_0_[1][40] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][410] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[410]),
        .Q(\shift_array_reg_n_0_[1][410] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][411] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[411]),
        .Q(\shift_array_reg_n_0_[1][411] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][412] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[412]),
        .Q(\shift_array_reg_n_0_[1][412] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][413] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[413]),
        .Q(\shift_array_reg_n_0_[1][413] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][414] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[414]),
        .Q(\shift_array_reg_n_0_[1][414] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][415] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[415]),
        .Q(\shift_array_reg_n_0_[1][415] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][416] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[416]),
        .Q(\shift_array_reg_n_0_[1][416] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][417] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[417]),
        .Q(\shift_array_reg_n_0_[1][417] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][418] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[418]),
        .Q(\shift_array_reg_n_0_[1][418] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][419] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[419]),
        .Q(\shift_array_reg_n_0_[1][419] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][41] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[41]),
        .Q(\shift_array_reg_n_0_[1][41] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][420] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[420]),
        .Q(\shift_array_reg_n_0_[1][420] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][421] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[421]),
        .Q(\shift_array_reg_n_0_[1][421] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][422] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[422]),
        .Q(\shift_array_reg_n_0_[1][422] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][423] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[423]),
        .Q(\shift_array_reg_n_0_[1][423] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][424] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[424]),
        .Q(\shift_array_reg_n_0_[1][424] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][425] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[425]),
        .Q(\shift_array_reg_n_0_[1][425] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][426] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[426]),
        .Q(\shift_array_reg_n_0_[1][426] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][427] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[427]),
        .Q(\shift_array_reg_n_0_[1][427] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][428] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[428]),
        .Q(\shift_array_reg_n_0_[1][428] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][429] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[429]),
        .Q(\shift_array_reg_n_0_[1][429] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][42] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[42]),
        .Q(\shift_array_reg_n_0_[1][42] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][430] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[430]),
        .Q(\shift_array_reg_n_0_[1][430] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][431] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[431]),
        .Q(\shift_array_reg_n_0_[1][431] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][432] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[432]),
        .Q(\shift_array_reg_n_0_[1][432] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][433] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[433]),
        .Q(\shift_array_reg_n_0_[1][433] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][434] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[434]),
        .Q(\shift_array_reg_n_0_[1][434] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][435] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[435]),
        .Q(\shift_array_reg_n_0_[1][435] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][436] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[436]),
        .Q(\shift_array_reg_n_0_[1][436] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][437] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[437]),
        .Q(\shift_array_reg_n_0_[1][437] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][438] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[438]),
        .Q(\shift_array_reg_n_0_[1][438] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][439] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[439]),
        .Q(\shift_array_reg_n_0_[1][439] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][43] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[43]),
        .Q(\shift_array_reg_n_0_[1][43] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][440] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[440]),
        .Q(\shift_array_reg_n_0_[1][440] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][441] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[441]),
        .Q(\shift_array_reg_n_0_[1][441] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][442] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[442]),
        .Q(\shift_array_reg_n_0_[1][442] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][443] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[443]),
        .Q(\shift_array_reg_n_0_[1][443] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][444] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[444]),
        .Q(\shift_array_reg_n_0_[1][444] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][445] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[445]),
        .Q(\shift_array_reg_n_0_[1][445] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][446] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[446]),
        .Q(\shift_array_reg_n_0_[1][446] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][447] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[447]),
        .Q(\shift_array_reg_n_0_[1][447] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][448] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[448]),
        .Q(\shift_array_reg_n_0_[1][448] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][449] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[449]),
        .Q(\shift_array_reg_n_0_[1][449] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][44] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[44]),
        .Q(\shift_array_reg_n_0_[1][44] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][450] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[450]),
        .Q(\shift_array_reg_n_0_[1][450] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][451] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[451]),
        .Q(\shift_array_reg_n_0_[1][451] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][452] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[452]),
        .Q(\shift_array_reg_n_0_[1][452] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][453] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[453]),
        .Q(\shift_array_reg_n_0_[1][453] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][454] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[454]),
        .Q(\shift_array_reg_n_0_[1][454] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][455] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[455]),
        .Q(\shift_array_reg_n_0_[1][455] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][456] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[456]),
        .Q(\shift_array_reg_n_0_[1][456] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][457] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[457]),
        .Q(\shift_array_reg_n_0_[1][457] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][458] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[458]),
        .Q(\shift_array_reg_n_0_[1][458] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][459] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[459]),
        .Q(\shift_array_reg_n_0_[1][459] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][45] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[45]),
        .Q(\shift_array_reg_n_0_[1][45] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][460] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[460]),
        .Q(\shift_array_reg_n_0_[1][460] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][461] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[461]),
        .Q(\shift_array_reg_n_0_[1][461] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][462] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[462]),
        .Q(\shift_array_reg_n_0_[1][462] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][463] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[463]),
        .Q(\shift_array_reg_n_0_[1][463] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][464] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[464]),
        .Q(\shift_array_reg_n_0_[1][464] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][465] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[465]),
        .Q(\shift_array_reg_n_0_[1][465] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][466] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[466]),
        .Q(\shift_array_reg_n_0_[1][466] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][467] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[467]),
        .Q(\shift_array_reg_n_0_[1][467] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][468] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[468]),
        .Q(\shift_array_reg_n_0_[1][468] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][469] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[469]),
        .Q(\shift_array_reg_n_0_[1][469] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][46] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[46]),
        .Q(\shift_array_reg_n_0_[1][46] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][470] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[470]),
        .Q(\shift_array_reg_n_0_[1][470] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][471] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[471]),
        .Q(\shift_array_reg_n_0_[1][471] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][472] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[472]),
        .Q(\shift_array_reg_n_0_[1][472] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][473] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[473]),
        .Q(\shift_array_reg_n_0_[1][473] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][474] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[474]),
        .Q(\shift_array_reg_n_0_[1][474] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][475] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[475]),
        .Q(\shift_array_reg_n_0_[1][475] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][476] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[476]),
        .Q(\shift_array_reg_n_0_[1][476] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][477] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[477]),
        .Q(\shift_array_reg_n_0_[1][477] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][478] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[478]),
        .Q(\shift_array_reg_n_0_[1][478] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][479] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[479]),
        .Q(\shift_array_reg_n_0_[1][479] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][47] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[47]),
        .Q(\shift_array_reg_n_0_[1][47] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][480] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[480]),
        .Q(\shift_array_reg_n_0_[1][480] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][481] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[481]),
        .Q(\shift_array_reg_n_0_[1][481] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][482] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[482]),
        .Q(\shift_array_reg_n_0_[1][482] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][483] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[483]),
        .Q(\shift_array_reg_n_0_[1][483] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][484] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[484]),
        .Q(\shift_array_reg_n_0_[1][484] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][485] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[485]),
        .Q(\shift_array_reg_n_0_[1][485] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][486] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[486]),
        .Q(\shift_array_reg_n_0_[1][486] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][487] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[487]),
        .Q(\shift_array_reg_n_0_[1][487] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][488] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[488]),
        .Q(\shift_array_reg_n_0_[1][488] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][489] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[489]),
        .Q(\shift_array_reg_n_0_[1][489] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][48] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[48]),
        .Q(\shift_array_reg_n_0_[1][48] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][490] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[490]),
        .Q(\shift_array_reg_n_0_[1][490] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][491] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[491]),
        .Q(\shift_array_reg_n_0_[1][491] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][492] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[492]),
        .Q(\shift_array_reg_n_0_[1][492] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][493] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[493]),
        .Q(\shift_array_reg_n_0_[1][493] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][494] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[494]),
        .Q(\shift_array_reg_n_0_[1][494] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][495] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[495]),
        .Q(\shift_array_reg_n_0_[1][495] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][496] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[496]),
        .Q(\shift_array_reg_n_0_[1][496] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][497] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[497]),
        .Q(\shift_array_reg_n_0_[1][497] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][498] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[498]),
        .Q(\shift_array_reg_n_0_[1][498] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][499] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[499]),
        .Q(\shift_array_reg_n_0_[1][499] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][49] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[49]),
        .Q(\shift_array_reg_n_0_[1][49] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[4]),
        .Q(\shift_array_reg_n_0_[1][4] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][500] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[500]),
        .Q(\shift_array_reg_n_0_[1][500] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][501] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[501]),
        .Q(\shift_array_reg_n_0_[1][501] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][502] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[502]),
        .Q(\shift_array_reg_n_0_[1][502] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][503] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[503]),
        .Q(\shift_array_reg_n_0_[1][503] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][504] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[504]),
        .Q(\shift_array_reg_n_0_[1][504] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][505] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[505]),
        .Q(\shift_array_reg_n_0_[1][505] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][506] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[506]),
        .Q(\shift_array_reg_n_0_[1][506] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][507] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[507]),
        .Q(\shift_array_reg_n_0_[1][507] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][508] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[508]),
        .Q(\shift_array_reg_n_0_[1][508] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][509] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[509]),
        .Q(\shift_array_reg_n_0_[1][509] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][50] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[50]),
        .Q(\shift_array_reg_n_0_[1][50] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][510] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[510]),
        .Q(\shift_array_reg_n_0_[1][510] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][511] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[511]),
        .Q(\shift_array_reg_n_0_[1][511] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][512] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[512]),
        .Q(\shift_array_reg_n_0_[1][512] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][513] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[513]),
        .Q(\shift_array_reg_n_0_[1][513] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][514] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[514]),
        .Q(\shift_array_reg_n_0_[1][514] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][515] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[515]),
        .Q(\shift_array_reg_n_0_[1][515] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][516] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[516]),
        .Q(\shift_array_reg_n_0_[1][516] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][517] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[517]),
        .Q(\shift_array_reg_n_0_[1][517] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][518] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[518]),
        .Q(\shift_array_reg_n_0_[1][518] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][519] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[519]),
        .Q(\shift_array_reg_n_0_[1][519] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][51] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[51]),
        .Q(\shift_array_reg_n_0_[1][51] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][520] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[520]),
        .Q(\shift_array_reg_n_0_[1][520] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][521] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[521]),
        .Q(\shift_array_reg_n_0_[1][521] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][522] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[522]),
        .Q(\shift_array_reg_n_0_[1][522] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][523] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[523]),
        .Q(\shift_array_reg_n_0_[1][523] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][524] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[524]),
        .Q(\shift_array_reg_n_0_[1][524] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][525] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[525]),
        .Q(\shift_array_reg_n_0_[1][525] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][526] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[526]),
        .Q(\shift_array_reg_n_0_[1][526] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][527] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[527]),
        .Q(\shift_array_reg_n_0_[1][527] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][528] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[528]),
        .Q(\shift_array_reg_n_0_[1][528] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][529] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[529]),
        .Q(\shift_array_reg_n_0_[1][529] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][52] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[52]),
        .Q(\shift_array_reg_n_0_[1][52] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][530] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[530]),
        .Q(\shift_array_reg_n_0_[1][530] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][531] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[531]),
        .Q(\shift_array_reg_n_0_[1][531] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][532] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[532]),
        .Q(\shift_array_reg_n_0_[1][532] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][533] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[533]),
        .Q(\shift_array_reg_n_0_[1][533] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][534] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[534]),
        .Q(\shift_array_reg_n_0_[1][534] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][535] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[535]),
        .Q(\shift_array_reg_n_0_[1][535] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][536] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[536]),
        .Q(\shift_array_reg_n_0_[1][536] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][537] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[537]),
        .Q(\shift_array_reg_n_0_[1][537] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][538] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[538]),
        .Q(\shift_array_reg_n_0_[1][538] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][539] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[539]),
        .Q(\shift_array_reg_n_0_[1][539] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][53] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[53]),
        .Q(\shift_array_reg_n_0_[1][53] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][540] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[540]),
        .Q(\shift_array_reg_n_0_[1][540] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][541] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[541]),
        .Q(\shift_array_reg_n_0_[1][541] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][542] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[542]),
        .Q(\shift_array_reg_n_0_[1][542] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][543] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[543]),
        .Q(\shift_array_reg_n_0_[1][543] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][544] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[544]),
        .Q(\shift_array_reg_n_0_[1][544] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][545] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[545]),
        .Q(\shift_array_reg_n_0_[1][545] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][546] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[546]),
        .Q(\shift_array_reg_n_0_[1][546] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][547] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[547]),
        .Q(\shift_array_reg_n_0_[1][547] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][548] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[548]),
        .Q(\shift_array_reg_n_0_[1][548] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][549] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[549]),
        .Q(\shift_array_reg_n_0_[1][549] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][54] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[54]),
        .Q(\shift_array_reg_n_0_[1][54] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][550] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[550]),
        .Q(\shift_array_reg_n_0_[1][550] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][551] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[551]),
        .Q(\shift_array_reg_n_0_[1][551] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][552] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[552]),
        .Q(\shift_array_reg_n_0_[1][552] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][553] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[553]),
        .Q(\shift_array_reg_n_0_[1][553] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][554] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[554]),
        .Q(\shift_array_reg_n_0_[1][554] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][555] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[555]),
        .Q(\shift_array_reg_n_0_[1][555] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][556] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[556]),
        .Q(\shift_array_reg_n_0_[1][556] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][557] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[557]),
        .Q(\shift_array_reg_n_0_[1][557] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][558] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[558]),
        .Q(\shift_array_reg_n_0_[1][558] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][559] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[559]),
        .Q(\shift_array_reg_n_0_[1][559] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][55] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[55]),
        .Q(\shift_array_reg_n_0_[1][55] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][560] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[560]),
        .Q(\shift_array_reg_n_0_[1][560] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][561] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[561]),
        .Q(\shift_array_reg_n_0_[1][561] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][562] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[562]),
        .Q(\shift_array_reg_n_0_[1][562] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][563] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[563]),
        .Q(\shift_array_reg_n_0_[1][563] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][564] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[564]),
        .Q(\shift_array_reg_n_0_[1][564] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][565] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[565]),
        .Q(\shift_array_reg_n_0_[1][565] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][566] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[566]),
        .Q(\shift_array_reg_n_0_[1][566] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][567] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[567]),
        .Q(\shift_array_reg_n_0_[1][567] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][568] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[568]),
        .Q(\shift_array_reg_n_0_[1][568] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][569] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[569]),
        .Q(\shift_array_reg_n_0_[1][569] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][56] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[56]),
        .Q(\shift_array_reg_n_0_[1][56] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][570] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[570]),
        .Q(\shift_array_reg_n_0_[1][570] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][571] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[571]),
        .Q(\shift_array_reg_n_0_[1][571] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][572] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[572]),
        .Q(\shift_array_reg_n_0_[1][572] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][573] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[573]),
        .Q(\shift_array_reg_n_0_[1][573] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][574] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[574]),
        .Q(\shift_array_reg_n_0_[1][574] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][575] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[575]),
        .Q(\shift_array_reg_n_0_[1][575] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][576] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[576]),
        .Q(\shift_array_reg_n_0_[1][576] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][577] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[577]),
        .Q(\shift_array_reg_n_0_[1][577] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][578] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[578]),
        .Q(\shift_array_reg_n_0_[1][578] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][579] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[579]),
        .Q(\shift_array_reg_n_0_[1][579] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][57] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[57]),
        .Q(\shift_array_reg_n_0_[1][57] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][580] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[580]),
        .Q(\shift_array_reg_n_0_[1][580] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][581] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[581]),
        .Q(\shift_array_reg_n_0_[1][581] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][582] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[582]),
        .Q(\shift_array_reg_n_0_[1][582] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][583] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[583]),
        .Q(\shift_array_reg_n_0_[1][583] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][584] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[584]),
        .Q(\shift_array_reg_n_0_[1][584] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][585] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[585]),
        .Q(\shift_array_reg_n_0_[1][585] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][586] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[586]),
        .Q(\shift_array_reg_n_0_[1][586] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][587] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[587]),
        .Q(\shift_array_reg_n_0_[1][587] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][588] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[588]),
        .Q(\shift_array_reg_n_0_[1][588] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][589] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[589]),
        .Q(\shift_array_reg_n_0_[1][589] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][58] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[58]),
        .Q(\shift_array_reg_n_0_[1][58] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][590] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[590]),
        .Q(\shift_array_reg_n_0_[1][590] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][591] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[591]),
        .Q(\shift_array_reg_n_0_[1][591] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][592] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[592]),
        .Q(\shift_array_reg_n_0_[1][592] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][593] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[593]),
        .Q(\shift_array_reg_n_0_[1][593] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][594] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[594]),
        .Q(\shift_array_reg_n_0_[1][594] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][595] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[595]),
        .Q(\shift_array_reg_n_0_[1][595] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][596] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[596]),
        .Q(\shift_array_reg_n_0_[1][596] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][597] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[597]),
        .Q(\shift_array_reg_n_0_[1][597] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][598] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[598]),
        .Q(\shift_array_reg_n_0_[1][598] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][599] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[599]),
        .Q(\shift_array_reg_n_0_[1][599] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][59] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[59]),
        .Q(\shift_array_reg_n_0_[1][59] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[5]),
        .Q(\shift_array_reg_n_0_[1][5] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][600] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[600]),
        .Q(\shift_array_reg_n_0_[1][600] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][601] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[601]),
        .Q(\shift_array_reg_n_0_[1][601] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][602] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[602]),
        .Q(\shift_array_reg_n_0_[1][602] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][603] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[603]),
        .Q(\shift_array_reg_n_0_[1][603] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][604] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[604]),
        .Q(\shift_array_reg_n_0_[1][604] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][605] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[605]),
        .Q(\shift_array_reg_n_0_[1][605] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][606] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[606]),
        .Q(\shift_array_reg_n_0_[1][606] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][607] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[607]),
        .Q(\shift_array_reg_n_0_[1][607] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][608] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[608]),
        .Q(\shift_array_reg_n_0_[1][608] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][609] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[609]),
        .Q(\shift_array_reg_n_0_[1][609] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][60] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[60]),
        .Q(\shift_array_reg_n_0_[1][60] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][610] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[610]),
        .Q(\shift_array_reg_n_0_[1][610] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][611] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[611]),
        .Q(\shift_array_reg_n_0_[1][611] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][612] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[612]),
        .Q(\shift_array_reg_n_0_[1][612] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][613] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[613]),
        .Q(\shift_array_reg_n_0_[1][613] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][614] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[614]),
        .Q(\shift_array_reg_n_0_[1][614] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][615] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[615]),
        .Q(\shift_array_reg_n_0_[1][615] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][616] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[616]),
        .Q(\shift_array_reg_n_0_[1][616] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][617] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[617]),
        .Q(\shift_array_reg_n_0_[1][617] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][618] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[618]),
        .Q(\shift_array_reg_n_0_[1][618] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][619] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[619]),
        .Q(\shift_array_reg_n_0_[1][619] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][61] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[61]),
        .Q(\shift_array_reg_n_0_[1][61] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][620] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[620]),
        .Q(\shift_array_reg_n_0_[1][620] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][621] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[621]),
        .Q(\shift_array_reg_n_0_[1][621] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][622] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[622]),
        .Q(\shift_array_reg_n_0_[1][622] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][623] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[623]),
        .Q(\shift_array_reg_n_0_[1][623] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][624] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[624]),
        .Q(\shift_array_reg_n_0_[1][624] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][625] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[625]),
        .Q(\shift_array_reg_n_0_[1][625] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][626] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[626]),
        .Q(\shift_array_reg_n_0_[1][626] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][627] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[627]),
        .Q(\shift_array_reg_n_0_[1][627] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][628] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[628]),
        .Q(\shift_array_reg_n_0_[1][628] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][629] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[629]),
        .Q(\shift_array_reg_n_0_[1][629] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][62] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[62]),
        .Q(\shift_array_reg_n_0_[1][62] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][630] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[630]),
        .Q(\shift_array_reg_n_0_[1][630] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][631] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[631]),
        .Q(\shift_array_reg_n_0_[1][631] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][632] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[632]),
        .Q(\shift_array_reg_n_0_[1][632] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][633] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[633]),
        .Q(\shift_array_reg_n_0_[1][633] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][634] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[634]),
        .Q(\shift_array_reg_n_0_[1][634] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][635] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[635]),
        .Q(\shift_array_reg_n_0_[1][635] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][636] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[636]),
        .Q(\shift_array_reg_n_0_[1][636] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][637] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[637]),
        .Q(\shift_array_reg_n_0_[1][637] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][638] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[638]),
        .Q(\shift_array_reg_n_0_[1][638] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][639] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[639]),
        .Q(\shift_array_reg_n_0_[1][639] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][63] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[63]),
        .Q(\shift_array_reg_n_0_[1][63] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][640] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[640]),
        .Q(\shift_array_reg_n_0_[1][640] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][641] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[641]),
        .Q(\shift_array_reg_n_0_[1][641] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][642] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[642]),
        .Q(\shift_array_reg_n_0_[1][642] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][643] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[643]),
        .Q(\shift_array_reg_n_0_[1][643] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][644] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[644]),
        .Q(\shift_array_reg_n_0_[1][644] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][645] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[645]),
        .Q(\shift_array_reg_n_0_[1][645] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][646] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[646]),
        .Q(\shift_array_reg_n_0_[1][646] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][647] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[647]),
        .Q(\shift_array_reg_n_0_[1][647] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][648] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[648]),
        .Q(\shift_array_reg_n_0_[1][648] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][649] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[649]),
        .Q(\shift_array_reg_n_0_[1][649] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][64] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[64]),
        .Q(\shift_array_reg_n_0_[1][64] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][650] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[650]),
        .Q(\shift_array_reg_n_0_[1][650] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][651] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[651]),
        .Q(\shift_array_reg_n_0_[1][651] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][652] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[652]),
        .Q(\shift_array_reg_n_0_[1][652] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][653] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[653]),
        .Q(\shift_array_reg_n_0_[1][653] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][654] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[654]),
        .Q(\shift_array_reg_n_0_[1][654] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][655] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[655]),
        .Q(\shift_array_reg_n_0_[1][655] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][656] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[656]),
        .Q(\shift_array_reg_n_0_[1][656] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][657] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[657]),
        .Q(\shift_array_reg_n_0_[1][657] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][658] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[658]),
        .Q(\shift_array_reg_n_0_[1][658] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][659] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[659]),
        .Q(\shift_array_reg_n_0_[1][659] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][65] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[65]),
        .Q(\shift_array_reg_n_0_[1][65] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][660] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[660]),
        .Q(\shift_array_reg_n_0_[1][660] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][661] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[661]),
        .Q(\shift_array_reg_n_0_[1][661] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][662] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[662]),
        .Q(\shift_array_reg_n_0_[1][662] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][663] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[663]),
        .Q(\shift_array_reg_n_0_[1][663] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][664] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[664]),
        .Q(\shift_array_reg_n_0_[1][664] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][665] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[665]),
        .Q(\shift_array_reg_n_0_[1][665] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][666] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[666]),
        .Q(\shift_array_reg_n_0_[1][666] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][667] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[667]),
        .Q(\shift_array_reg_n_0_[1][667] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][668] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[668]),
        .Q(\shift_array_reg_n_0_[1][668] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][669] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[669]),
        .Q(\shift_array_reg_n_0_[1][669] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][66] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[66]),
        .Q(\shift_array_reg_n_0_[1][66] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][670] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[670]),
        .Q(\shift_array_reg_n_0_[1][670] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][671] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[671]),
        .Q(\shift_array_reg_n_0_[1][671] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][672] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[672]),
        .Q(\shift_array_reg_n_0_[1][672] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][673] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[673]),
        .Q(\shift_array_reg_n_0_[1][673] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][674] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[674]),
        .Q(\shift_array_reg_n_0_[1][674] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][675] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[675]),
        .Q(\shift_array_reg_n_0_[1][675] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][676] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[676]),
        .Q(\shift_array_reg_n_0_[1][676] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][677] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[677]),
        .Q(\shift_array_reg_n_0_[1][677] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][678] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[678]),
        .Q(\shift_array_reg_n_0_[1][678] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][679] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[679]),
        .Q(\shift_array_reg_n_0_[1][679] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][67] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[67]),
        .Q(\shift_array_reg_n_0_[1][67] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][680] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[680]),
        .Q(\shift_array_reg_n_0_[1][680] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][681] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[681]),
        .Q(\shift_array_reg_n_0_[1][681] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][682] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[682]),
        .Q(\shift_array_reg_n_0_[1][682] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][683] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[683]),
        .Q(\shift_array_reg_n_0_[1][683] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][684] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[684]),
        .Q(\shift_array_reg_n_0_[1][684] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][685] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[685]),
        .Q(\shift_array_reg_n_0_[1][685] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][686] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[686]),
        .Q(\shift_array_reg_n_0_[1][686] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][687] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[687]),
        .Q(\shift_array_reg_n_0_[1][687] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][688] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[688]),
        .Q(\shift_array_reg_n_0_[1][688] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][689] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[689]),
        .Q(\shift_array_reg_n_0_[1][689] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][68] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[68]),
        .Q(\shift_array_reg_n_0_[1][68] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][690] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[690]),
        .Q(\shift_array_reg_n_0_[1][690] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][691] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[691]),
        .Q(\shift_array_reg_n_0_[1][691] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][692] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[692]),
        .Q(\shift_array_reg_n_0_[1][692] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][693] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[693]),
        .Q(\shift_array_reg_n_0_[1][693] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][694] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[694]),
        .Q(\shift_array_reg_n_0_[1][694] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][695] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[695]),
        .Q(\shift_array_reg_n_0_[1][695] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][696] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[696]),
        .Q(\shift_array_reg_n_0_[1][696] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][697] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[697]),
        .Q(\shift_array_reg_n_0_[1][697] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][698] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[698]),
        .Q(\shift_array_reg_n_0_[1][698] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][699] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[699]),
        .Q(\shift_array_reg_n_0_[1][699] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][69] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[69]),
        .Q(\shift_array_reg_n_0_[1][69] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[6]),
        .Q(\shift_array_reg_n_0_[1][6] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][700] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[700]),
        .Q(\shift_array_reg_n_0_[1][700] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][701] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[701]),
        .Q(\shift_array_reg_n_0_[1][701] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][702] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[702]),
        .Q(\shift_array_reg_n_0_[1][702] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][703] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[703]),
        .Q(\shift_array_reg_n_0_[1][703] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][704] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[704]),
        .Q(\shift_array_reg_n_0_[1][704] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][705] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[705]),
        .Q(\shift_array_reg_n_0_[1][705] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][706] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[706]),
        .Q(\shift_array_reg_n_0_[1][706] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][707] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[707]),
        .Q(\shift_array_reg_n_0_[1][707] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][708] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[708]),
        .Q(\shift_array_reg_n_0_[1][708] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][709] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[709]),
        .Q(\shift_array_reg_n_0_[1][709] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][70] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[70]),
        .Q(\shift_array_reg_n_0_[1][70] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][710] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[710]),
        .Q(\shift_array_reg_n_0_[1][710] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][711] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[711]),
        .Q(\shift_array_reg_n_0_[1][711] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][712] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[712]),
        .Q(\shift_array_reg_n_0_[1][712] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][713] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[713]),
        .Q(\shift_array_reg_n_0_[1][713] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][714] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[714]),
        .Q(\shift_array_reg_n_0_[1][714] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][715] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[715]),
        .Q(\shift_array_reg_n_0_[1][715] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][716] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[716]),
        .Q(\shift_array_reg_n_0_[1][716] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][717] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[717]),
        .Q(\shift_array_reg_n_0_[1][717] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][718] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[718]),
        .Q(\shift_array_reg_n_0_[1][718] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][719] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[719]),
        .Q(\shift_array_reg_n_0_[1][719] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][71] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[71]),
        .Q(\shift_array_reg_n_0_[1][71] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][720] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[720]),
        .Q(\shift_array_reg_n_0_[1][720] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][721] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[721]),
        .Q(\shift_array_reg_n_0_[1][721] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][722] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[722]),
        .Q(\shift_array_reg_n_0_[1][722] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][723] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[723]),
        .Q(\shift_array_reg_n_0_[1][723] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][724] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[724]),
        .Q(\shift_array_reg_n_0_[1][724] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][725] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[725]),
        .Q(\shift_array_reg_n_0_[1][725] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][726] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[726]),
        .Q(\shift_array_reg_n_0_[1][726] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][727] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[727]),
        .Q(\shift_array_reg_n_0_[1][727] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][728] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[728]),
        .Q(\shift_array_reg_n_0_[1][728] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][729] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[729]),
        .Q(\shift_array_reg_n_0_[1][729] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][72] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[72]),
        .Q(\shift_array_reg_n_0_[1][72] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][730] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[730]),
        .Q(\shift_array_reg_n_0_[1][730] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][731] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[731]),
        .Q(\shift_array_reg_n_0_[1][731] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][732] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[732]),
        .Q(\shift_array_reg_n_0_[1][732] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][733] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[733]),
        .Q(\shift_array_reg_n_0_[1][733] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][734] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[734]),
        .Q(\shift_array_reg_n_0_[1][734] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][735] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[735]),
        .Q(\shift_array_reg_n_0_[1][735] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][736] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[736]),
        .Q(\shift_array_reg_n_0_[1][736] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][737] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[737]),
        .Q(\shift_array_reg_n_0_[1][737] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][738] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[738]),
        .Q(\shift_array_reg_n_0_[1][738] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][739] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[739]),
        .Q(\shift_array_reg_n_0_[1][739] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][73] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[73]),
        .Q(\shift_array_reg_n_0_[1][73] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][740] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[740]),
        .Q(\shift_array_reg_n_0_[1][740] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][741] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[741]),
        .Q(\shift_array_reg_n_0_[1][741] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][742] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[742]),
        .Q(\shift_array_reg_n_0_[1][742] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][743] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[743]),
        .Q(\shift_array_reg_n_0_[1][743] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][744] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[744]),
        .Q(\shift_array_reg_n_0_[1][744] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][745] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[745]),
        .Q(\shift_array_reg_n_0_[1][745] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][746] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[746]),
        .Q(\shift_array_reg_n_0_[1][746] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][747] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[747]),
        .Q(\shift_array_reg_n_0_[1][747] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][748] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[748]),
        .Q(\shift_array_reg_n_0_[1][748] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][749] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[749]),
        .Q(\shift_array_reg_n_0_[1][749] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][74] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[74]),
        .Q(\shift_array_reg_n_0_[1][74] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][750] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[750]),
        .Q(\shift_array_reg_n_0_[1][750] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][751] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[751]),
        .Q(\shift_array_reg_n_0_[1][751] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][752] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[752]),
        .Q(\shift_array_reg_n_0_[1][752] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][753] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[753]),
        .Q(\shift_array_reg_n_0_[1][753] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][754] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[754]),
        .Q(\shift_array_reg_n_0_[1][754] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][755] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[755]),
        .Q(\shift_array_reg_n_0_[1][755] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][756] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[756]),
        .Q(\shift_array_reg_n_0_[1][756] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][757] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[757]),
        .Q(\shift_array_reg_n_0_[1][757] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][758] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[758]),
        .Q(\shift_array_reg_n_0_[1][758] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][759] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[759]),
        .Q(\shift_array_reg_n_0_[1][759] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][75] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[75]),
        .Q(\shift_array_reg_n_0_[1][75] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][760] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[760]),
        .Q(\shift_array_reg_n_0_[1][760] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][761] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[761]),
        .Q(\shift_array_reg_n_0_[1][761] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][762] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[762]),
        .Q(\shift_array_reg_n_0_[1][762] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][763] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[763]),
        .Q(\shift_array_reg_n_0_[1][763] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][764] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[764]),
        .Q(\shift_array_reg_n_0_[1][764] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][765] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[765]),
        .Q(\shift_array_reg_n_0_[1][765] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][766] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[766]),
        .Q(\shift_array_reg_n_0_[1][766] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][767] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[767]),
        .Q(\shift_array_reg_n_0_[1][767] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][768] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[768]),
        .Q(\shift_array_reg_n_0_[1][768] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][769] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[769]),
        .Q(\shift_array_reg_n_0_[1][769] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][76] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[76]),
        .Q(\shift_array_reg_n_0_[1][76] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][770] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[770]),
        .Q(\shift_array_reg_n_0_[1][770] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][771] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[771]),
        .Q(\shift_array_reg_n_0_[1][771] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][772] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[772]),
        .Q(\shift_array_reg_n_0_[1][772] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][773] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[773]),
        .Q(\shift_array_reg_n_0_[1][773] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][774] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[774]),
        .Q(\shift_array_reg_n_0_[1][774] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][775] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[775]),
        .Q(\shift_array_reg_n_0_[1][775] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][776] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[776]),
        .Q(\shift_array_reg_n_0_[1][776] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][777] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[777]),
        .Q(\shift_array_reg_n_0_[1][777] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][778] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[778]),
        .Q(\shift_array_reg_n_0_[1][778] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][779] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[779]),
        .Q(\shift_array_reg_n_0_[1][779] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][77] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[77]),
        .Q(\shift_array_reg_n_0_[1][77] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][780] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[780]),
        .Q(\shift_array_reg_n_0_[1][780] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][781] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[781]),
        .Q(\shift_array_reg_n_0_[1][781] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][782] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[782]),
        .Q(\shift_array_reg_n_0_[1][782] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][783] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[783]),
        .Q(\shift_array_reg_n_0_[1][783] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][784] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[784]),
        .Q(\shift_array_reg_n_0_[1][784] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][785] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[785]),
        .Q(\shift_array_reg_n_0_[1][785] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][786] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[786]),
        .Q(\shift_array_reg_n_0_[1][786] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][787] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[787]),
        .Q(\shift_array_reg_n_0_[1][787] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][788] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[788]),
        .Q(\shift_array_reg_n_0_[1][788] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][789] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[789]),
        .Q(\shift_array_reg_n_0_[1][789] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][78] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[78]),
        .Q(\shift_array_reg_n_0_[1][78] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][790] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[790]),
        .Q(\shift_array_reg_n_0_[1][790] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][791] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[791]),
        .Q(\shift_array_reg_n_0_[1][791] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][792] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[792]),
        .Q(\shift_array_reg_n_0_[1][792] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][793] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[793]),
        .Q(\shift_array_reg_n_0_[1][793] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][794] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[794]),
        .Q(\shift_array_reg_n_0_[1][794] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][795] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[795]),
        .Q(\shift_array_reg_n_0_[1][795] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][796] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[796]),
        .Q(\shift_array_reg_n_0_[1][796] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][797] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[797]),
        .Q(\shift_array_reg_n_0_[1][797] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][798] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[798]),
        .Q(\shift_array_reg_n_0_[1][798] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][799] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[799]),
        .Q(\shift_array_reg_n_0_[1][799] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][79] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[79]),
        .Q(\shift_array_reg_n_0_[1][79] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[7]),
        .Q(\shift_array_reg_n_0_[1][7] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][800] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[800]),
        .Q(\shift_array_reg_n_0_[1][800] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][801] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[801]),
        .Q(\shift_array_reg_n_0_[1][801] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][802] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[802]),
        .Q(\shift_array_reg_n_0_[1][802] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][803] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[803]),
        .Q(\shift_array_reg_n_0_[1][803] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][804] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[804]),
        .Q(\shift_array_reg_n_0_[1][804] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][805] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[805]),
        .Q(\shift_array_reg_n_0_[1][805] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][806] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[806]),
        .Q(\shift_array_reg_n_0_[1][806] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][807] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[807]),
        .Q(\shift_array_reg_n_0_[1][807] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][808] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[808]),
        .Q(\shift_array_reg_n_0_[1][808] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][809] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[809]),
        .Q(\shift_array_reg_n_0_[1][809] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][80] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[80]),
        .Q(\shift_array_reg_n_0_[1][80] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][810] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[810]),
        .Q(\shift_array_reg_n_0_[1][810] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][811] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[811]),
        .Q(\shift_array_reg_n_0_[1][811] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][812] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[812]),
        .Q(\shift_array_reg_n_0_[1][812] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][813] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[813]),
        .Q(\shift_array_reg_n_0_[1][813] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][814] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[814]),
        .Q(\shift_array_reg_n_0_[1][814] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][815] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[815]),
        .Q(\shift_array_reg_n_0_[1][815] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][816] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[816]),
        .Q(\shift_array_reg_n_0_[1][816] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][817] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[817]),
        .Q(\shift_array_reg_n_0_[1][817] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][818] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[818]),
        .Q(\shift_array_reg_n_0_[1][818] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][819] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[819]),
        .Q(\shift_array_reg_n_0_[1][819] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][81] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[81]),
        .Q(\shift_array_reg_n_0_[1][81] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][820] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[820]),
        .Q(\shift_array_reg_n_0_[1][820] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][821] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[821]),
        .Q(\shift_array_reg_n_0_[1][821] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][822] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[822]),
        .Q(\shift_array_reg_n_0_[1][822] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][823] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[823]),
        .Q(\shift_array_reg_n_0_[1][823] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][824] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[824]),
        .Q(\shift_array_reg_n_0_[1][824] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][825] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[825]),
        .Q(\shift_array_reg_n_0_[1][825] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][826] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[826]),
        .Q(\shift_array_reg_n_0_[1][826] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][827] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[827]),
        .Q(\shift_array_reg_n_0_[1][827] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][828] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[828]),
        .Q(\shift_array_reg_n_0_[1][828] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][829] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[829]),
        .Q(\shift_array_reg_n_0_[1][829] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][82] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[82]),
        .Q(\shift_array_reg_n_0_[1][82] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][830] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[830]),
        .Q(\shift_array_reg_n_0_[1][830] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][831] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[831]),
        .Q(\shift_array_reg_n_0_[1][831] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][832] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[832]),
        .Q(\shift_array_reg_n_0_[1][832] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][833] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[833]),
        .Q(\shift_array_reg_n_0_[1][833] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][834] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[834]),
        .Q(\shift_array_reg_n_0_[1][834] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][835] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[835]),
        .Q(\shift_array_reg_n_0_[1][835] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][836] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[836]),
        .Q(\shift_array_reg_n_0_[1][836] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][837] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[837]),
        .Q(\shift_array_reg_n_0_[1][837] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][838] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[838]),
        .Q(\shift_array_reg_n_0_[1][838] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][839] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[839]),
        .Q(\shift_array_reg_n_0_[1][839] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][83] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[83]),
        .Q(\shift_array_reg_n_0_[1][83] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][840] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[840]),
        .Q(\shift_array_reg_n_0_[1][840] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][841] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[841]),
        .Q(\shift_array_reg_n_0_[1][841] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][842] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[842]),
        .Q(\shift_array_reg_n_0_[1][842] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][843] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[843]),
        .Q(\shift_array_reg_n_0_[1][843] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][844] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[844]),
        .Q(\shift_array_reg_n_0_[1][844] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][845] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[845]),
        .Q(\shift_array_reg_n_0_[1][845] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][846] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[846]),
        .Q(\shift_array_reg_n_0_[1][846] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][847] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[847]),
        .Q(\shift_array_reg_n_0_[1][847] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][848] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[848]),
        .Q(\shift_array_reg_n_0_[1][848] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][849] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[849]),
        .Q(\shift_array_reg_n_0_[1][849] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][84] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[84]),
        .Q(\shift_array_reg_n_0_[1][84] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][850] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[850]),
        .Q(\shift_array_reg_n_0_[1][850] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][851] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[851]),
        .Q(\shift_array_reg_n_0_[1][851] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][852] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[852]),
        .Q(\shift_array_reg_n_0_[1][852] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][853] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[853]),
        .Q(\shift_array_reg_n_0_[1][853] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][854] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[854]),
        .Q(\shift_array_reg_n_0_[1][854] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][855] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[855]),
        .Q(\shift_array_reg_n_0_[1][855] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][856] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[856]),
        .Q(\shift_array_reg_n_0_[1][856] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][857] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[857]),
        .Q(\shift_array_reg_n_0_[1][857] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][858] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[858]),
        .Q(\shift_array_reg_n_0_[1][858] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][859] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[859]),
        .Q(\shift_array_reg_n_0_[1][859] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][85] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[85]),
        .Q(\shift_array_reg_n_0_[1][85] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][860] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[860]),
        .Q(\shift_array_reg_n_0_[1][860] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][861] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[861]),
        .Q(\shift_array_reg_n_0_[1][861] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][862] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[862]),
        .Q(\shift_array_reg_n_0_[1][862] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][863] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[863]),
        .Q(\shift_array_reg_n_0_[1][863] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][864] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[864]),
        .Q(\shift_array_reg_n_0_[1][864] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][865] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[865]),
        .Q(\shift_array_reg_n_0_[1][865] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][866] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[866]),
        .Q(\shift_array_reg_n_0_[1][866] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][867] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[867]),
        .Q(\shift_array_reg_n_0_[1][867] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][868] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[868]),
        .Q(\shift_array_reg_n_0_[1][868] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][869] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[869]),
        .Q(\shift_array_reg_n_0_[1][869] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][86] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[86]),
        .Q(\shift_array_reg_n_0_[1][86] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][870] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[870]),
        .Q(\shift_array_reg_n_0_[1][870] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][871] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[871]),
        .Q(\shift_array_reg_n_0_[1][871] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][872] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[872]),
        .Q(\shift_array_reg_n_0_[1][872] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][873] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[873]),
        .Q(\shift_array_reg_n_0_[1][873] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][874] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[874]),
        .Q(\shift_array_reg_n_0_[1][874] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][875] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[875]),
        .Q(\shift_array_reg_n_0_[1][875] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][876] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[876]),
        .Q(\shift_array_reg_n_0_[1][876] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][877] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[877]),
        .Q(\shift_array_reg_n_0_[1][877] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][878] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[878]),
        .Q(\shift_array_reg_n_0_[1][878] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][879] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[879]),
        .Q(\shift_array_reg_n_0_[1][879] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][87] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[87]),
        .Q(\shift_array_reg_n_0_[1][87] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][880] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[880]),
        .Q(\shift_array_reg_n_0_[1][880] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][881] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[881]),
        .Q(\shift_array_reg_n_0_[1][881] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][882] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[882]),
        .Q(\shift_array_reg_n_0_[1][882] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][883] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[883]),
        .Q(\shift_array_reg_n_0_[1][883] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][884] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[884]),
        .Q(\shift_array_reg_n_0_[1][884] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][885] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[885]),
        .Q(\shift_array_reg_n_0_[1][885] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][886] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[886]),
        .Q(\shift_array_reg_n_0_[1][886] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][887] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[887]),
        .Q(\shift_array_reg_n_0_[1][887] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][888] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[888]),
        .Q(\shift_array_reg_n_0_[1][888] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][889] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[889]),
        .Q(\shift_array_reg_n_0_[1][889] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][88] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[88]),
        .Q(\shift_array_reg_n_0_[1][88] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][890] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[890]),
        .Q(\shift_array_reg_n_0_[1][890] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][891] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[891]),
        .Q(\shift_array_reg_n_0_[1][891] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][892] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[892]),
        .Q(\shift_array_reg_n_0_[1][892] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][893] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[893]),
        .Q(\shift_array_reg_n_0_[1][893] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][894] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[894]),
        .Q(\shift_array_reg_n_0_[1][894] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][895] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[895]),
        .Q(\shift_array_reg_n_0_[1][895] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][896] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[896]),
        .Q(\shift_array_reg_n_0_[1][896] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][897] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[897]),
        .Q(\shift_array_reg_n_0_[1][897] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][898] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[898]),
        .Q(\shift_array_reg_n_0_[1][898] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][899] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[899]),
        .Q(\shift_array_reg_n_0_[1][899] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][89] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[89]),
        .Q(\shift_array_reg_n_0_[1][89] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[8]),
        .Q(\shift_array_reg_n_0_[1][8] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][900] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[900]),
        .Q(\shift_array_reg_n_0_[1][900] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][901] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[901]),
        .Q(\shift_array_reg_n_0_[1][901] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][902] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[902]),
        .Q(\shift_array_reg_n_0_[1][902] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][903] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[903]),
        .Q(\shift_array_reg_n_0_[1][903] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][904] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[904]),
        .Q(\shift_array_reg_n_0_[1][904] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][905] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[905]),
        .Q(\shift_array_reg_n_0_[1][905] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][906] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[906]),
        .Q(\shift_array_reg_n_0_[1][906] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][907] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[907]),
        .Q(\shift_array_reg_n_0_[1][907] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][908] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[908]),
        .Q(\shift_array_reg_n_0_[1][908] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][909] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[909]),
        .Q(\shift_array_reg_n_0_[1][909] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][90] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[90]),
        .Q(\shift_array_reg_n_0_[1][90] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][910] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[910]),
        .Q(\shift_array_reg_n_0_[1][910] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][911] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[911]),
        .Q(\shift_array_reg_n_0_[1][911] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][912] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[912]),
        .Q(\shift_array_reg_n_0_[1][912] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][913] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[913]),
        .Q(\shift_array_reg_n_0_[1][913] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][914] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[914]),
        .Q(\shift_array_reg_n_0_[1][914] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][915] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[915]),
        .Q(\shift_array_reg_n_0_[1][915] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][916] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[916]),
        .Q(\shift_array_reg_n_0_[1][916] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][917] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[917]),
        .Q(\shift_array_reg_n_0_[1][917] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][918] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[918]),
        .Q(\shift_array_reg_n_0_[1][918] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][919] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[919]),
        .Q(\shift_array_reg_n_0_[1][919] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][91] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[91]),
        .Q(\shift_array_reg_n_0_[1][91] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][920] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[920]),
        .Q(\shift_array_reg_n_0_[1][920] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][921] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[921]),
        .Q(\shift_array_reg_n_0_[1][921] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][922] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[922]),
        .Q(\shift_array_reg_n_0_[1][922] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][923] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[923]),
        .Q(\shift_array_reg_n_0_[1][923] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][924] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[924]),
        .Q(\shift_array_reg_n_0_[1][924] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][925] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[925]),
        .Q(\shift_array_reg_n_0_[1][925] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][926] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[926]),
        .Q(\shift_array_reg_n_0_[1][926] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][927] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[927]),
        .Q(\shift_array_reg_n_0_[1][927] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][928] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[928]),
        .Q(\shift_array_reg_n_0_[1][928] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][929] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[929]),
        .Q(\shift_array_reg_n_0_[1][929] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][92] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[92]),
        .Q(\shift_array_reg_n_0_[1][92] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][930] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[930]),
        .Q(\shift_array_reg_n_0_[1][930] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][931] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[931]),
        .Q(\shift_array_reg_n_0_[1][931] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][932] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[932]),
        .Q(\shift_array_reg_n_0_[1][932] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][933] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[933]),
        .Q(\shift_array_reg_n_0_[1][933] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][934] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[934]),
        .Q(\shift_array_reg_n_0_[1][934] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][935] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[935]),
        .Q(\shift_array_reg_n_0_[1][935] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][936] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[936]),
        .Q(\shift_array_reg_n_0_[1][936] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][937] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[937]),
        .Q(\shift_array_reg_n_0_[1][937] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][938] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[938]),
        .Q(\shift_array_reg_n_0_[1][938] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][939] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[939]),
        .Q(\shift_array_reg_n_0_[1][939] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][93] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[93]),
        .Q(\shift_array_reg_n_0_[1][93] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][940] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[940]),
        .Q(\shift_array_reg_n_0_[1][940] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][941] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[941]),
        .Q(\shift_array_reg_n_0_[1][941] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][942] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[942]),
        .Q(\shift_array_reg_n_0_[1][942] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][943] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[943]),
        .Q(\shift_array_reg_n_0_[1][943] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][944] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[944]),
        .Q(\shift_array_reg_n_0_[1][944] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][945] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[945]),
        .Q(\shift_array_reg_n_0_[1][945] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][946] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[946]),
        .Q(\shift_array_reg_n_0_[1][946] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][947] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[947]),
        .Q(\shift_array_reg_n_0_[1][947] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][948] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[948]),
        .Q(\shift_array_reg_n_0_[1][948] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][949] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[949]),
        .Q(\shift_array_reg_n_0_[1][949] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][94] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[94]),
        .Q(\shift_array_reg_n_0_[1][94] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][950] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[950]),
        .Q(\shift_array_reg_n_0_[1][950] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][951] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[951]),
        .Q(\shift_array_reg_n_0_[1][951] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][952] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[952]),
        .Q(\shift_array_reg_n_0_[1][952] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][953] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[953]),
        .Q(\shift_array_reg_n_0_[1][953] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][954] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[954]),
        .Q(\shift_array_reg_n_0_[1][954] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][955] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[955]),
        .Q(\shift_array_reg_n_0_[1][955] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][956] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[956]),
        .Q(\shift_array_reg_n_0_[1][956] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][957] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[957]),
        .Q(\shift_array_reg_n_0_[1][957] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][958] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[958]),
        .Q(\shift_array_reg_n_0_[1][958] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][959] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[959]),
        .Q(\shift_array_reg_n_0_[1][959] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][95] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[95]),
        .Q(\shift_array_reg_n_0_[1][95] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][960] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[960]),
        .Q(\shift_array_reg_n_0_[1][960] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][961] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[961]),
        .Q(\shift_array_reg_n_0_[1][961] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][962] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[962]),
        .Q(\shift_array_reg_n_0_[1][962] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][963] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[963]),
        .Q(\shift_array_reg_n_0_[1][963] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][964] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[964]),
        .Q(\shift_array_reg_n_0_[1][964] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][965] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[965]),
        .Q(\shift_array_reg_n_0_[1][965] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][966] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[966]),
        .Q(\shift_array_reg_n_0_[1][966] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][967] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[967]),
        .Q(\shift_array_reg_n_0_[1][967] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][968] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[968]),
        .Q(\shift_array_reg_n_0_[1][968] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][969] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[969]),
        .Q(\shift_array_reg_n_0_[1][969] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][96] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[96]),
        .Q(\shift_array_reg_n_0_[1][96] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][970] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[970]),
        .Q(\shift_array_reg_n_0_[1][970] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][971] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[971]),
        .Q(\shift_array_reg_n_0_[1][971] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][972] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[972]),
        .Q(\shift_array_reg_n_0_[1][972] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][973] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[973]),
        .Q(\shift_array_reg_n_0_[1][973] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][974] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[974]),
        .Q(\shift_array_reg_n_0_[1][974] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][975] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[975]),
        .Q(\shift_array_reg_n_0_[1][975] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][976] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[976]),
        .Q(\shift_array_reg_n_0_[1][976] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][977] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[977]),
        .Q(\shift_array_reg_n_0_[1][977] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][978] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[978]),
        .Q(\shift_array_reg_n_0_[1][978] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][979] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[979]),
        .Q(\shift_array_reg_n_0_[1][979] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][97] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[97]),
        .Q(\shift_array_reg_n_0_[1][97] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][980] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[980]),
        .Q(\shift_array_reg_n_0_[1][980] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][981] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[981]),
        .Q(\shift_array_reg_n_0_[1][981] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][982] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[982]),
        .Q(\shift_array_reg_n_0_[1][982] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][983] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[983]),
        .Q(\shift_array_reg_n_0_[1][983] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][984] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[984]),
        .Q(\shift_array_reg_n_0_[1][984] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][985] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[985]),
        .Q(\shift_array_reg_n_0_[1][985] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][986] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[986]),
        .Q(\shift_array_reg_n_0_[1][986] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][987] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[987]),
        .Q(\shift_array_reg_n_0_[1][987] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][988] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[988]),
        .Q(\shift_array_reg_n_0_[1][988] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][989] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[989]),
        .Q(\shift_array_reg_n_0_[1][989] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][98] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[98]),
        .Q(\shift_array_reg_n_0_[1][98] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][990] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[990]),
        .Q(\shift_array_reg_n_0_[1][990] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][991] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[991]),
        .Q(\shift_array_reg_n_0_[1][991] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][992] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[992]),
        .Q(\shift_array_reg_n_0_[1][992] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][993] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[993]),
        .Q(\shift_array_reg_n_0_[1][993] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][994] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[994]),
        .Q(\shift_array_reg_n_0_[1][994] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][995] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[995]),
        .Q(\shift_array_reg_n_0_[1][995] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][996] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[996]),
        .Q(\shift_array_reg_n_0_[1][996] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][997] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[997]),
        .Q(\shift_array_reg_n_0_[1][997] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][998] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[998]),
        .Q(\shift_array_reg_n_0_[1][998] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][999] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[999]),
        .Q(\shift_array_reg_n_0_[1][999] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][99] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[99]),
        .Q(\shift_array_reg_n_0_[1][99] ),
        .R(\<const0> ));
  (* SHREG_EXTRACT = "yes" *) 
  FDRE #(
    .INIT(1'b0)) 
    \shift_array_reg[1][9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_point_i[9]),
        .Q(\shift_array_reg_n_0_[1][9] ),
        .R(\<const0> ));
endmodule

(* ADDR_WIDTH_A = "15" *) (* ADDR_WIDTH_B = "15" *) (* AUTO_SLEEP_TIME = "0" *) 
(* BYTE_WRITE_WIDTH_A = "1" *) (* BYTE_WRITE_WIDTH_B = "1" *) (* CASCADE_HEIGHT = "0" *) 
(* CLOCKING_MODE = "0" *) (* CORE_GENERATION_INFO = "xpm_memory_base,xpm_memory_base,{MEMORY_TYPE=2,MEMORY_SIZE=32768,MEMORY_PRIMITIVE=2,CLOCKING_MODE=0,ECC_MODE=0,ECC_TYPE=NONE,ECC_BIT_RANGE=[7:0],MEMORY_INIT_PARAM=,IGNORE_INIT_SYNTH=0,USE_MEM_INIT_MMI=0,USE_MEM_INIT=1,MEMORY_OPTIMIZATION=true,WAKEUP_TIME=0,AUTO_SLEEP_TIME=0,MESSAGE_CONTROL=0,VERSION=0,USE_EMBEDDED_CONSTRAINT=0,CASCADE_HEIGHT=0,SIM_ASSERT_CHK=0,WRITE_PROTECT=1,RAM_DECOMP=auto,WRITE_DATA_WIDTH_A=1,READ_DATA_WIDTH_A=1,BYTE_WRITE_WIDTH_A=1,ADDR_WIDTH_A=15,READ_RESET_VALUE_A=0,READ_LATENCY_A=3,WRITE_MODE_A=1,RST_MODE_A=SYNC,WRITE_DATA_WIDTH_B=1,READ_DATA_WIDTH_B=1,BYTE_WRITE_WIDTH_B=1,ADDR_WIDTH_B=15,READ_RESET_VALUE_B=0,READ_LATENCY_B=3,WRITE_MODE_B=1,RST_MODE_B=SYNC,P_MEMORY_PRIMITIVE=block,P_MIN_WIDTH_DATA_A=1,P_MIN_WIDTH_DATA_B=1,P_MIN_WIDTH_DATA=1,P_MIN_WIDTH_DATA_ECC=1,P_MAX_DEPTH_DATA=32768,P_ECC_MODE=no_ecc,P_MEMORY_OPT=yes,P_WIDTH_COL_WRITE_A=1,P_WIDTH_COL_WRITE_B=1,P_NUM_COLS_WRITE_A=1,P_NUM_COLS_WRITE_B=1,P_NUM_ROWS_WRITE_A=1,P_NUM_ROWS_WRITE_B=1,P_NUM_ROWS_READ_A=1,P_NUM_ROWS_READ_B=1,P_WIDTH_ADDR_WRITE_A=15,P_WIDTH_ADDR_WRITE_B=15,P_WIDTH_ADDR_READ_A=15,P_WIDTH_ADDR_READ_B=15,P_WIDTH_ADDR_LSB_WRITE_A=0,P_WIDTH_ADDR_LSB_WRITE_B=0,P_WIDTH_ADDR_LSB_READ_A=0,P_WIDTH_ADDR_LSB_READ_B=0,P_ENABLE_BYTE_WRITE_A=0,P_ENABLE_BYTE_WRITE_B=0,P_SDP_WRITE_MODE=yes,rsta_loop_iter=4,rstb_loop_iter=4,NUM_CHAR_LOC=0,MAX_NUM_CHAR=0,P_MIN_WIDTH_DATA_SHFT=5,P_MIN_WIDTH_DATA_LDW=1}" *) (* ECC_BIT_RANGE = "[7:0]" *) 
(* ECC_MODE = "0" *) (* ECC_TYPE = "NONE" *) (* IGNORE_INIT_SYNTH = "0" *) 
(* MAX_NUM_CHAR = "0" *) (* MEMORY_INIT_FILE = "none" *) (* MEMORY_INIT_PARAM = "" *) 
(* MEMORY_OPTIMIZATION = "true" *) (* MEMORY_PRIMITIVE = "2" *) (* MEMORY_SIZE = "32768" *) 
(* MEMORY_TYPE = "2" *) (* MESSAGE_CONTROL = "0" *) (* NUM_CHAR_LOC = "0" *) 
(* ORIG_REF_NAME = "xpm_memory_base" *) (* P_ECC_MODE = "0" *) (* P_ENABLE_BYTE_WRITE_A = "0" *) 
(* P_ENABLE_BYTE_WRITE_B = "0" *) (* P_MAX_DEPTH_DATA = "32768" *) (* P_MEMORY_OPT = "yes" *) 
(* P_MEMORY_PRIMITIVE = "0" *) (* P_MIN_WIDTH_DATA = "1" *) (* P_MIN_WIDTH_DATA_A = "1" *) 
(* P_MIN_WIDTH_DATA_B = "1" *) (* P_MIN_WIDTH_DATA_ECC = "1" *) (* P_MIN_WIDTH_DATA_LDW = "1" *) 
(* P_MIN_WIDTH_DATA_SHFT = "5" *) (* P_NUM_COLS_WRITE_A = "1" *) (* P_NUM_COLS_WRITE_B = "1" *) 
(* P_NUM_ROWS_READ_A = "1" *) (* P_NUM_ROWS_READ_B = "1" *) (* P_NUM_ROWS_WRITE_A = "1" *) 
(* P_NUM_ROWS_WRITE_B = "1" *) (* P_SDP_WRITE_MODE = "yes" *) (* P_WIDTH_ADDR_LSB_READ_A = "0" *) 
(* P_WIDTH_ADDR_LSB_READ_B = "0" *) (* P_WIDTH_ADDR_LSB_WRITE_A = "0" *) (* P_WIDTH_ADDR_LSB_WRITE_B = "0" *) 
(* P_WIDTH_ADDR_READ_A = "15" *) (* P_WIDTH_ADDR_READ_B = "15" *) (* P_WIDTH_ADDR_WRITE_A = "15" *) 
(* P_WIDTH_ADDR_WRITE_B = "15" *) (* P_WIDTH_COL_WRITE_A = "1" *) (* P_WIDTH_COL_WRITE_B = "1" *) 
(* RAM_DECOMP = "auto" *) (* READ_DATA_WIDTH_A = "1" *) (* READ_DATA_WIDTH_B = "1" *) 
(* READ_LATENCY_A = "3" *) (* READ_LATENCY_B = "3" *) (* READ_RESET_VALUE_A = "0" *) 
(* READ_RESET_VALUE_B = "0" *) (* RST_MODE_A = "SYNC" *) (* RST_MODE_B = "SYNC" *) 
(* SIM_ASSERT_CHK = "0" *) (* USE_EMBEDDED_CONSTRAINT = "0" *) (* USE_MEM_INIT = "1" *) 
(* USE_MEM_INIT_MMI = "0" *) (* VERSION = "0" *) (* WAKEUP_TIME = "0" *) 
(* WRITE_DATA_WIDTH_A = "1" *) (* WRITE_DATA_WIDTH_B = "1" *) (* WRITE_MODE_A = "1" *) 
(* WRITE_MODE_B = "1" *) (* WRITE_PROTECT = "1" *) (* XPM_MODULE = "TRUE" *) 
(* keep_hierarchy = "soft" *) (* rsta_loop_iter = "4" *) (* rstb_loop_iter = "4" *) 
module ponos_xpm_memory_base
   (sleep,
    clka,
    rsta,
    ena,
    regcea,
    wea,
    addra,
    dina,
    injectsbiterra,
    injectdbiterra,
    douta,
    sbiterra,
    dbiterra,
    clkb,
    rstb,
    enb,
    regceb,
    web,
    addrb,
    dinb,
    injectsbiterrb,
    injectdbiterrb,
    doutb,
    sbiterrb,
    dbiterrb);
  input sleep;
  input clka;
  input rsta;
  input ena;
  input regcea;
  input [0:0]wea;
  input [14:0]addra;
  input [0:0]dina;
  input injectsbiterra;
  input injectdbiterra;
  output [0:0]douta;
  output sbiterra;
  output dbiterra;
  input clkb;
  input rstb;
  input enb;
  input regceb;
  input [0:0]web;
  input [14:0]addrb;
  input [0:0]dinb;
  input injectsbiterrb;
  input injectdbiterrb;
  output [0:0]doutb;
  output sbiterrb;
  output dbiterrb;

  wire \<const0> ;
  wire \<const1> ;
  wire VCC_2;
  wire [14:0]addra;
  wire [14:0]addrb;
  wire clka;
  wire [0:0]dina;
  wire [0:0]douta;
  wire \gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe[1][0]_i_1_n_0 ;
  wire \gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[0] ;
  wire \gen_wr_a.gen_word_narrow.mem_reg_bram_0_n_99 ;
  wire rsta;
  wire sleep;
  wire [0:0]wea;
  wire [0:0]web;

  assign dbiterra = \<const0> ;
  assign dbiterrb = \<const0> ;
  assign doutb[0] = \<const0> ;
  assign sbiterra = \<const0> ;
  assign sbiterrb = \<const0> ;
  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  VCC VCC_1
       (.P(VCC_2));
  LUT2 #(
    .INIT(4'h2)) 
    \gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe[1][0]_i_1 
       (.I0(\gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[0] ),
        .I1(rsta),
        .O(\gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe[1][0]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[1][0] 
       (.C(clka),
        .CE(\<const1> ),
        .D(\gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe[1][0]_i_1_n_0 ),
        .Q(douta),
        .R(\<const0> ));
  (* \MEM.PORTA.ADDRESS_BEGIN  = "0" *) 
  (* \MEM.PORTA.ADDRESS_END  = "32767" *) 
  (* \MEM.PORTA.DATA_BIT_LAYOUT  = "p0_d1" *) 
  (* \MEM.PORTA.DATA_LSB  = "0" *) 
  (* \MEM.PORTA.DATA_MSB  = "0" *) 
  (* \MEM.PORTB.ADDRESS_BEGIN  = "0" *) 
  (* \MEM.PORTB.ADDRESS_END  = "32767" *) 
  (* \MEM.PORTB.DATA_BIT_LAYOUT  = "p0_d1" *) 
  (* \MEM.PORTB.DATA_LSB  = "0" *) 
  (* \MEM.PORTB.DATA_MSB  = "0" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-7 {cell *THIS*}}" *) 
  (* RDADDR_COLLISION_HWCONFIG = "DELAYED_WRITE" *) 
  (* RTL_RAM_BITS = "32768" *) 
  (* RTL_RAM_NAME = "i_tdpram_flag_mem/xpm_memory_base_inst/gen_wr_a.gen_word_narrow.mem_reg_bram_0" *) 
  (* RTL_RAM_TYPE = "RAM_TDP" *) 
  (* ram_addr_begin = "0" *) 
  (* ram_addr_end = "32767" *) 
  (* ram_offset = "0" *) 
  (* ram_slice_begin = "0" *) 
  (* ram_slice_end = "0" *) 
  RAMB36E2 #(
    .CASCADE_ORDER_A("NONE"),
    .CASCADE_ORDER_B("NONE"),
    .CLOCK_DOMAINS("COMMON"),
    .DOA_REG(0),
    .DOB_REG(1),
    .ENADDRENA("FALSE"),
    .ENADDRENB("FALSE"),
    .EN_ECC_PIPE("FALSE"),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .INIT_FILE("NONE"),
    .RDADDRCHANGEA("FALSE"),
    .RDADDRCHANGEB("FALSE"),
    .READ_WIDTH_A(1),
    .READ_WIDTH_B(1),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SLEEP_ASYNC("FALSE"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("READ_FIRST"),
    .WRITE_WIDTH_A(1),
    .WRITE_WIDTH_B(1)) 
    \gen_wr_a.gen_word_narrow.mem_reg_bram_0 
       (.ADDRARDADDR(addrb),
        .ADDRBWRADDR(addra),
        .ADDRENA(\<const1> ),
        .ADDRENB(\<const1> ),
        .CASDIMUXA(\<const0> ),
        .CASDIMUXB(\<const0> ),
        .CASDINA({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .CASDINB({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .CASDINPA({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .CASDINPB({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .CASDOMUXA(\<const0> ),
        .CASDOMUXB(\<const0> ),
        .CASDOMUXEN_A(\<const1> ),
        .CASDOMUXEN_B(\<const1> ),
        .CASINDBITERR(\<const0> ),
        .CASINSBITERR(\<const0> ),
        .CASOREGIMUXA(\<const0> ),
        .CASOREGIMUXB(\<const0> ),
        .CASOREGIMUXEN_A(\<const1> ),
        .CASOREGIMUXEN_B(\<const1> ),
        .CLKARDCLK(clka),
        .CLKBWRCLK(clka),
        .DINADIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .DINBDIN({\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,\<const0> ,dina}),
        .DINPADINP({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .DINPBDINP({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .DOUTADOUT(\gen_wr_a.gen_word_narrow.mem_reg_bram_0_n_99 ),
        .DOUTBDOUT(\gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[0] ),
        .ECCPIPECE(VCC_2),
        .ENARDEN(\<const1> ),
        .ENBWREN(\<const1> ),
        .INJECTDBITERR(\<const0> ),
        .INJECTSBITERR(\<const0> ),
        .REGCEAREGCE(\<const1> ),
        .REGCEB(\<const1> ),
        .RSTRAMARSTRAM(\<const0> ),
        .RSTRAMB(\<const0> ),
        .RSTREGARSTREG(\<const0> ),
        .RSTREGB(\<const0> ),
        .SLEEP(\<const0> ),
        .WEA({web,web,web,web}),
        .WEBWE({\<const0> ,\<const0> ,\<const0> ,\<const0> ,wea,wea,wea,wea}));
endmodule

(* ADDR_WIDTH_A = "15" *) (* ADDR_WIDTH_B = "15" *) (* AUTO_SLEEP_TIME = "0" *) 
(* BYTE_WRITE_WIDTH_A = "1" *) (* BYTE_WRITE_WIDTH_B = "1" *) (* CASCADE_HEIGHT = "0" *) 
(* CLOCKING_MODE = "common_clock" *) (* CORE_GENERATION_INFO = "xpm_memory_tdpram,xpm_memory_tdpram,{MEMORY_SIZE=32768,MEMORY_PRIMITIVE=block,CLOCKING_MODE=common_clock,ECC_MODE=no_ecc,ECC_TYPE=NONE,ECC_BIT_RANGE=[7:0],MEMORY_INIT_PARAM=,USE_MEM_INIT=1,USE_MEM_INIT_MMI=0,WAKEUP_TIME=disable_sleep,AUTO_SLEEP_TIME=0,MESSAGE_CONTROL=0,USE_EMBEDDED_CONSTRAINT=0,MEMORY_OPTIMIZATION=true,CASCADE_HEIGHT=0,RAM_DECOMP=auto,SIM_ASSERT_CHK=0,WRITE_PROTECT=1,IGNORE_INIT_SYNTH=0,WRITE_DATA_WIDTH_A=1,READ_DATA_WIDTH_A=1,BYTE_WRITE_WIDTH_A=1,ADDR_WIDTH_A=15,READ_RESET_VALUE_A=0,READ_LATENCY_A=3,WRITE_MODE_A=read_first,RST_MODE_A=SYNC,WRITE_DATA_WIDTH_B=1,READ_DATA_WIDTH_B=1,BYTE_WRITE_WIDTH_B=1,ADDR_WIDTH_B=15,READ_RESET_VALUE_B=0,READ_LATENCY_B=3,WRITE_MODE_B=read_first,RST_MODE_B=SYNC,P_MEMORY_PRIMITIVE=2,P_CLOCKING_MODE=0,P_ECC_MODE=0,P_WAKEUP_TIME=0,P_WRITE_MODE_A=1,P_WRITE_MODE_B=1,P_MEMORY_OPTIMIZATION=1}" *) (* ECC_BIT_RANGE = "[7:0]" *) 
(* ECC_MODE = "no_ecc" *) (* ECC_TYPE = "NONE" *) (* IGNORE_INIT_SYNTH = "0" *) 
(* MEMORY_INIT_FILE = "none" *) (* MEMORY_INIT_PARAM = "" *) (* MEMORY_OPTIMIZATION = "true" *) 
(* MEMORY_PRIMITIVE = "block" *) (* MEMORY_SIZE = "32768" *) (* MESSAGE_CONTROL = "0" *) 
(* ORIG_REF_NAME = "xpm_memory_tdpram" *) (* P_CLOCKING_MODE = "0" *) (* P_ECC_MODE = "0" *) 
(* P_MEMORY_OPTIMIZATION = "1" *) (* P_MEMORY_PRIMITIVE = "2" *) (* P_WAKEUP_TIME = "0" *) 
(* P_WRITE_MODE_A = "1" *) (* P_WRITE_MODE_B = "1" *) (* RAM_DECOMP = "auto" *) 
(* READ_DATA_WIDTH_A = "1" *) (* READ_DATA_WIDTH_B = "1" *) (* READ_LATENCY_A = "3" *) 
(* READ_LATENCY_B = "3" *) (* READ_RESET_VALUE_A = "0" *) (* READ_RESET_VALUE_B = "0" *) 
(* RST_MODE_A = "SYNC" *) (* RST_MODE_B = "SYNC" *) (* SIM_ASSERT_CHK = "0" *) 
(* USE_EMBEDDED_CONSTRAINT = "0" *) (* USE_MEM_INIT = "1" *) (* USE_MEM_INIT_MMI = "0" *) 
(* WAKEUP_TIME = "disable_sleep" *) (* WRITE_DATA_WIDTH_A = "1" *) (* WRITE_DATA_WIDTH_B = "1" *) 
(* WRITE_MODE_A = "read_first" *) (* WRITE_MODE_B = "read_first" *) (* WRITE_PROTECT = "1" *) 
(* XPM_MODULE = "TRUE" *) 
module ponos_xpm_memory_tdpram
   (sleep,
    clka,
    rsta,
    ena,
    regcea,
    wea,
    addra,
    dina,
    injectsbiterra,
    injectdbiterra,
    douta,
    sbiterra,
    dbiterra,
    clkb,
    rstb,
    enb,
    regceb,
    web,
    addrb,
    dinb,
    injectsbiterrb,
    injectdbiterrb,
    doutb,
    sbiterrb,
    dbiterrb);
  input sleep;
  input clka;
  input rsta;
  input ena;
  input regcea;
  input [0:0]wea;
  input [14:0]addra;
  input [0:0]dina;
  input injectsbiterra;
  input injectdbiterra;
  output [0:0]douta;
  output sbiterra;
  output dbiterra;
  input clkb;
  input rstb;
  input enb;
  input regceb;
  input [0:0]web;
  input [14:0]addrb;
  input [0:0]dinb;
  input injectsbiterrb;
  input injectdbiterrb;
  output [0:0]doutb;
  output sbiterrb;
  output dbiterrb;

  wire \<const0> ;
  wire \<const1> ;
  wire [14:0]addra;
  wire [14:0]addrb;
  wire clka;
  wire [0:0]dina;
  wire [0:0]douta;
  wire rsta;
  wire sleep;
  wire [0:0]wea;
  wire [0:0]web;

  assign dbiterra = \<const0> ;
  assign dbiterrb = \<const0> ;
  assign doutb[0] = \<const0> ;
  assign sbiterra = \<const0> ;
  assign sbiterrb = \<const0> ;
  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* ADDR_WIDTH_A = "15" *) 
  (* ADDR_WIDTH_B = "15" *) 
  (* AUTO_SLEEP_TIME = "0" *) 
  (* BYTE_WRITE_WIDTH_A = "1" *) 
  (* BYTE_WRITE_WIDTH_B = "1" *) 
  (* CASCADE_HEIGHT = "0" *) 
  (* CLOCKING_MODE = "0" *) 
  (* ECC_BIT_RANGE = "[7:0]" *) 
  (* ECC_MODE = "0" *) 
  (* ECC_TYPE = "NONE" *) 
  (* IGNORE_INIT_SYNTH = "0" *) 
  (* KEEP_HIERARCHY = "soft" *) 
  (* MAX_NUM_CHAR = "0" *) 
  (* \MEM.ADDRESS_SPACE  *) 
  (* \MEM.ADDRESS_SPACE_BEGIN  = "0" *) 
  (* \MEM.ADDRESS_SPACE_DATA_LSB  = "0" *) 
  (* \MEM.ADDRESS_SPACE_DATA_MSB  = "0" *) 
  (* \MEM.ADDRESS_SPACE_END  = "32767" *) 
  (* \MEM.CORE_MEMORY_WIDTH  = "1" *) 
  (* MEMORY_INIT_FILE = "none" *) 
  (* MEMORY_INIT_PARAM = "" *) 
  (* MEMORY_OPTIMIZATION = "true" *) 
  (* MEMORY_PRIMITIVE = "2" *) 
  (* MEMORY_SIZE = "32768" *) 
  (* MEMORY_TYPE = "2" *) 
  (* MESSAGE_CONTROL = "0" *) 
  (* NUM_CHAR_LOC = "0" *) 
  (* P_ECC_MODE = "no_ecc" *) 
  (* P_ENABLE_BYTE_WRITE_A = "0" *) 
  (* P_ENABLE_BYTE_WRITE_B = "0" *) 
  (* P_MAX_DEPTH_DATA = "32768" *) 
  (* P_MEMORY_OPT = "yes" *) 
  (* P_MEMORY_PRIMITIVE = "block" *) 
  (* P_MIN_WIDTH_DATA = "1" *) 
  (* P_MIN_WIDTH_DATA_A = "1" *) 
  (* P_MIN_WIDTH_DATA_B = "1" *) 
  (* P_MIN_WIDTH_DATA_ECC = "1" *) 
  (* P_MIN_WIDTH_DATA_LDW = "1" *) 
  (* P_MIN_WIDTH_DATA_SHFT = "5" *) 
  (* P_NUM_COLS_WRITE_A = "1" *) 
  (* P_NUM_COLS_WRITE_B = "1" *) 
  (* P_NUM_ROWS_READ_A = "1" *) 
  (* P_NUM_ROWS_READ_B = "1" *) 
  (* P_NUM_ROWS_WRITE_A = "1" *) 
  (* P_NUM_ROWS_WRITE_B = "1" *) 
  (* P_SDP_WRITE_MODE = "yes" *) 
  (* P_WIDTH_ADDR_LSB_READ_A = "0" *) 
  (* P_WIDTH_ADDR_LSB_READ_B = "0" *) 
  (* P_WIDTH_ADDR_LSB_WRITE_A = "0" *) 
  (* P_WIDTH_ADDR_LSB_WRITE_B = "0" *) 
  (* P_WIDTH_ADDR_READ_A = "15" *) 
  (* P_WIDTH_ADDR_READ_B = "15" *) 
  (* P_WIDTH_ADDR_WRITE_A = "15" *) 
  (* P_WIDTH_ADDR_WRITE_B = "15" *) 
  (* P_WIDTH_COL_WRITE_A = "1" *) 
  (* P_WIDTH_COL_WRITE_B = "1" *) 
  (* RAM_DECOMP = "auto" *) 
  (* READ_DATA_WIDTH_A = "1" *) 
  (* READ_DATA_WIDTH_B = "1" *) 
  (* READ_LATENCY_A = "3" *) 
  (* READ_LATENCY_B = "3" *) 
  (* READ_RESET_VALUE_A = "0" *) 
  (* READ_RESET_VALUE_B = "0" *) 
  (* RST_MODE_A = "SYNC" *) 
  (* RST_MODE_B = "SYNC" *) 
  (* SIM_ASSERT_CHK = "0" *) 
  (* USE_EMBEDDED_CONSTRAINT = "0" *) 
  (* USE_MEM_INIT = "1" *) 
  (* USE_MEM_INIT_MMI = "0" *) 
  (* VERSION = "0" *) 
  (* WAKEUP_TIME = "0" *) 
  (* WRITE_DATA_WIDTH_A = "1" *) 
  (* WRITE_DATA_WIDTH_B = "1" *) 
  (* WRITE_MODE_A = "1" *) 
  (* WRITE_MODE_B = "1" *) 
  (* WRITE_PROTECT = "1" *) 
  (* XPM_MODULE = "TRUE" *) 
  (* rsta_loop_iter = "4" *) 
  (* rstb_loop_iter = "4" *) 
  ponos_xpm_memory_base xpm_memory_base_inst
       (.addra(addra),
        .addrb(addrb),
        .clka(clka),
        .clkb(\<const0> ),
        .dina(dina),
        .dinb(\<const0> ),
        .douta(douta),
        .ena(\<const1> ),
        .enb(\<const1> ),
        .injectdbiterra(\<const0> ),
        .injectdbiterrb(\<const0> ),
        .injectsbiterra(\<const0> ),
        .injectsbiterrb(\<const0> ),
        .regcea(\<const1> ),
        .regceb(\<const0> ),
        .rsta(rsta),
        .rstb(\<const0> ),
        .sleep(sleep),
        .wea(wea),
        .web(web));
endmodule

(* LP_BUCKET_ADDR_WIDTH = "12" *) (* LP_BUCKET_SET_ADDR_WIDTH = "3" *) (* LP_DUMMY_INDEX_VAL = "3'b111" *) 
(* LP_FLAG_ADDR_WIDTH = "15" *) (* LP_FLAG_MEM_READ_LATENCY = "3" *) (* LP_VALID_DL_DEPTH = "4" *) 
(* P_DATA_PNT_W = "388" *) (* P_NUM_AFF_COORD = "3" *) (* P_NUM_WIN = "7" *) 
(* P_RED_SCLR_W = "13" *) 
(* STRUCTURAL_NETLIST = "yes" *)
module scheduler
   (clk,
    rst_n,
    prsi_point_i,
    prsi_red_scalar_i,
    prsi_index_i,
    prsi_valid_i,
    prsi_last_i,
    prsi_ready_o,
    accept_flags_o,
    accept_valid_o,
    acc_point_o,
    acc_bucket_addr_o,
    acc_bucket_set_addr_o,
    acc_add_sub_o,
    acc_valid_o,
    bm_bucket_addr_i,
    bm_bucket_set_addr_i,
    bm_valid_i,
    init_done_i);
  input clk;
  input rst_n;
  input [1163:0]prsi_point_i;
  input [12:0]prsi_red_scalar_i;
  input [2:0]prsi_index_i;
  input prsi_valid_i;
  input prsi_last_i;
  output prsi_ready_o;
  output [6:0]accept_flags_o;
  output accept_valid_o;
  output [1163:0]acc_point_o;
  output [11:0]acc_bucket_addr_o;
  output [2:0]acc_bucket_set_addr_o;
  output acc_add_sub_o;
  output acc_valid_o;
  input [11:0]bm_bucket_addr_i;
  input [2:0]bm_bucket_set_addr_i;
  input bm_valid_i;
  input init_done_i;

  wire \<const0> ;
  wire \<const1> ;
  wire \DELAY_BLOCK[3].shift_array_reg[4] ;
  wire acc_add_sub_o;
  wire [11:0]acc_bucket_addr_o;
  wire [2:0]acc_bucket_set_addr_o;
  wire [1163:0]acc_point_o;
  wire acc_valid_o;
  wire acc_valid_o0;
  wire [6:0]accept_flags_o;
  wire accept_valid_o;
  wire accept_valid_o0;
  wire [11:0]bm_bucket_addr_i;
  wire [2:0]bm_bucket_set_addr_i;
  wire bm_valid_i;
  wire [2:0]calc_bucket_set_addr_i_dld;
  wire calc_is_dummy_dld;
  wire calc_is_zero;
  wire calc_is_zero_dld;
  wire [14:0]clear_bucket_flag_addr;
  wire \clear_bucket_flag_addr[0]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[10]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[11]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[12]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[13]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[14]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[1]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[2]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[3]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[4]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[5]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[6]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[7]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[8]_i_1_n_0 ;
  wire \clear_bucket_flag_addr[9]_i_1_n_0 ;
  wire clear_bucket_flag_we;
  wire clk;
  wire [11:0]data0;
  wire i_shiftreg_calc_bucket_addr_n_0;
  wire i_shiftreg_calc_bucket_addr_n_1;
  wire i_shiftreg_calc_bucket_addr_n_10;
  wire i_shiftreg_calc_bucket_addr_n_11;
  wire i_shiftreg_calc_bucket_addr_n_13;
  wire i_shiftreg_calc_bucket_addr_n_2;
  wire i_shiftreg_calc_bucket_addr_n_3;
  wire i_shiftreg_calc_bucket_addr_n_4;
  wire i_shiftreg_calc_bucket_addr_n_5;
  wire i_shiftreg_calc_bucket_addr_n_6;
  wire i_shiftreg_calc_bucket_addr_n_7;
  wire i_shiftreg_calc_bucket_addr_n_8;
  wire i_shiftreg_calc_bucket_addr_n_9;
  wire i_shiftreg_calc_bucket_set_addr_n_3;
  wire i_shiftreg_calc_bucket_set_addr_n_4;
  wire i_shiftreg_calc_bucket_set_addr_n_5;
  wire i_shiftreg_calc_bucket_set_addr_n_6;
  wire i_shiftreg_calc_bucket_set_addr_n_7;
  wire i_shiftreg_calc_bucket_set_addr_n_8;
  wire i_shiftreg_calc_bucket_set_addr_n_9;
  wire i_shiftreg_calc_is_zero_n_1;
  wire i_shiftreg_calc_is_zero_n_2;
  wire i_shiftreg_calc_is_zero_n_3;
  wire i_shiftreg_calc_is_zero_n_4;
  wire i_shiftreg_calc_is_zero_n_5;
  wire init_done_i;
  wire \last_dld_reg_n_0_[0] ;
  wire \last_dld_reg_n_0_[1] ;
  wire \last_dld_reg_n_0_[2] ;
  wire \last_dld_reg_n_0_[3] ;
  wire [14:0]mark_check_bucket_flag_addr;
  wire \mark_check_bucket_flag_addr[11]_i_1_n_0 ;
  wire \mark_check_bucket_flag_addr[12]_i_1_n_0 ;
  wire \mark_check_bucket_flag_addr[13]_i_1_n_0 ;
  wire \mark_check_bucket_flag_addr[14]_i_1_n_0 ;
  wire mark_check_bucket_flag_out;
  wire mark_check_bucket_flag_we;
  wire mark_check_bucket_flag_we_i_10_n_0;
  wire mark_check_bucket_flag_we_i_11_n_0;
  wire mark_check_bucket_flag_we_i_1_n_0;
  wire mark_check_bucket_flag_we_i_2_n_0;
  wire mark_check_bucket_flag_we_i_3_n_0;
  wire mark_check_bucket_flag_we_i_4_n_0;
  wire mark_check_bucket_flag_we_i_5_n_0;
  wire mark_check_bucket_flag_we_i_6_n_0;
  wire mark_check_bucket_flag_we_i_7_n_0;
  wire mark_check_bucket_flag_we_i_8_n_0;
  wire mark_check_bucket_flag_we_i_9_n_0;
  wire p_7_in;
  wire processing_first_accept_flag;
  wire processing_first_accept_flag_i_1_n_0;
  wire [2:0]prsi_index_i;
  wire prsi_last_i;
  wire [1163:0]prsi_point_i;
  wire prsi_ready_o;
  wire prsi_ready_o_i_1_n_0;
  wire [12:0]prsi_red_scalar_i;
  wire prsi_valid_i;
  wire rst_n;
  wire \valid_dld_reg_n_0_[0] ;
  wire \valid_dld_reg_n_0_[1] ;
  wire \valid_dld_reg_n_0_[2] ;
  wire \valid_dld_reg_n_0_[3] ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  FDRE #(
    .INIT(1'b0)) 
    acc_add_sub_o_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(\DELAY_BLOCK[3].shift_array_reg[4] ),
        .Q(acc_add_sub_o),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_11),
        .Q(acc_bucket_addr_o[0]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_1),
        .Q(acc_bucket_addr_o[10]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_0),
        .Q(acc_bucket_addr_o[11]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_10),
        .Q(acc_bucket_addr_o[1]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_9),
        .Q(acc_bucket_addr_o[2]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_8),
        .Q(acc_bucket_addr_o[3]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_7),
        .Q(acc_bucket_addr_o[4]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_6),
        .Q(acc_bucket_addr_o[5]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_5),
        .Q(acc_bucket_addr_o[6]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_4),
        .Q(acc_bucket_addr_o[7]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_3),
        .Q(acc_bucket_addr_o[8]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_addr_o_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_addr_n_2),
        .Q(acc_bucket_addr_o[9]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_set_addr_o_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(calc_bucket_set_addr_i_dld[0]),
        .Q(acc_bucket_set_addr_o[0]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_set_addr_o_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(calc_bucket_set_addr_i_dld[1]),
        .Q(acc_bucket_set_addr_o[1]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \acc_bucket_set_addr_o_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(calc_bucket_set_addr_i_dld[2]),
        .Q(acc_bucket_set_addr_o[2]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    acc_valid_o_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(acc_valid_o0),
        .Q(acc_valid_o),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \accept_flags_o_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_set_addr_n_5),
        .Q(accept_flags_o[0]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \accept_flags_o_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_is_zero_n_5),
        .Q(accept_flags_o[1]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \accept_flags_o_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_set_addr_n_4),
        .Q(accept_flags_o[2]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \accept_flags_o_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_is_zero_n_4),
        .Q(accept_flags_o[3]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \accept_flags_o_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_is_zero_n_3),
        .Q(accept_flags_o[4]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \accept_flags_o_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_bucket_set_addr_n_3),
        .Q(accept_flags_o[5]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \accept_flags_o_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(i_shiftreg_calc_is_zero_n_1),
        .Q(accept_flags_o[6]),
        .R(prsi_ready_o_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    accept_valid_o_i_1
       (.I0(\valid_dld_reg_n_0_[3] ),
        .I1(\last_dld_reg_n_0_[3] ),
        .O(accept_valid_o0));
  FDRE #(
    .INIT(1'b0)) 
    accept_valid_o_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(accept_valid_o0),
        .Q(accept_valid_o),
        .R(prsi_ready_o_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[0]_i_1 
       (.I0(bm_bucket_addr_i[0]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[0]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[10]_i_1 
       (.I0(bm_bucket_addr_i[10]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[10]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[11]_i_1 
       (.I0(bm_bucket_addr_i[11]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[12]_i_1 
       (.I0(bm_bucket_set_addr_i[0]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[13]_i_1 
       (.I0(bm_bucket_set_addr_i[1]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[14]_i_1 
       (.I0(bm_bucket_set_addr_i[2]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[14]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[1]_i_1 
       (.I0(bm_bucket_addr_i[1]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[1]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[2]_i_1 
       (.I0(bm_bucket_addr_i[2]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[2]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[3]_i_1 
       (.I0(bm_bucket_addr_i[3]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[3]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[4]_i_1 
       (.I0(bm_bucket_addr_i[4]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[4]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[5]_i_1 
       (.I0(bm_bucket_addr_i[5]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[5]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[6]_i_1 
       (.I0(bm_bucket_addr_i[6]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[6]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[7]_i_1 
       (.I0(bm_bucket_addr_i[7]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[7]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[8]_i_1 
       (.I0(bm_bucket_addr_i[8]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[8]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \clear_bucket_flag_addr[9]_i_1 
       (.I0(bm_bucket_addr_i[9]),
        .I1(bm_valid_i),
        .O(\clear_bucket_flag_addr[9]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[0]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[0]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[10]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[10]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[11]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[11]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[12]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[12]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[13]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[13]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[14]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[14]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[1]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[1]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[2]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[2]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[3]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[3]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[4]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[4]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[5]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[5]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[6]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[6]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[7]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[7]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[8]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[8]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \clear_bucket_flag_addr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\clear_bucket_flag_addr[9]_i_1_n_0 ),
        .Q(clear_bucket_flag_addr[9]),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    clear_bucket_flag_we_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(bm_valid_i),
        .Q(clear_bucket_flag_we),
        .R(prsi_ready_o_i_1_n_0));
  ponos_shiftreg i_shiftreg_calc_add_sub
       (.\DELAY_BLOCK[3].shift_array_reg[4] (\DELAY_BLOCK[3].shift_array_reg[4] ),
        .clk(clk),
        .prsi_red_scalar_i(prsi_red_scalar_i[12]));
  ponos_shiftreg__parameterized0 i_shiftreg_calc_bucket_addr
       (.D({i_shiftreg_calc_bucket_addr_n_0,i_shiftreg_calc_bucket_addr_n_1,i_shiftreg_calc_bucket_addr_n_2,i_shiftreg_calc_bucket_addr_n_3,i_shiftreg_calc_bucket_addr_n_4,i_shiftreg_calc_bucket_addr_n_5,i_shiftreg_calc_bucket_addr_n_6,i_shiftreg_calc_bucket_addr_n_7,i_shiftreg_calc_bucket_addr_n_8,i_shiftreg_calc_bucket_addr_n_9,i_shiftreg_calc_bucket_addr_n_10,i_shiftreg_calc_bucket_addr_n_11}),
        .calc_is_zero(calc_is_zero),
        .clk(clk),
        .data0(data0),
        .prsi_red_scalar_i(prsi_red_scalar_i),
        .prsi_red_scalar_i_4_sp_1(i_shiftreg_calc_bucket_addr_n_13));
  ponos_shiftreg__parameterized1 i_shiftreg_calc_bucket_set_addr
       (.\DELAY_BLOCK[3].shift_array_reg[4][0]_0 (i_shiftreg_calc_bucket_set_addr_n_6),
        .\DELAY_BLOCK[3].shift_array_reg[4][0]_1 (i_shiftreg_calc_bucket_set_addr_n_9),
        .\DELAY_BLOCK[3].shift_array_reg[4][1]_0 (i_shiftreg_calc_bucket_set_addr_n_4),
        .\DELAY_BLOCK[3].shift_array_reg[4][1]_1 (i_shiftreg_calc_bucket_set_addr_n_5),
        .\DELAY_BLOCK[3].shift_array_reg[4][2]_0 (i_shiftreg_calc_bucket_set_addr_n_7),
        .\DELAY_BLOCK[3].shift_array_reg[4][2]_1 (i_shiftreg_calc_bucket_set_addr_n_8),
        .Q(\valid_dld_reg_n_0_[3] ),
        .accept_flags_o({accept_flags_o[5],accept_flags_o[2],accept_flags_o[0]}),
        .\accept_flags_o_reg[2] (i_shiftreg_calc_is_zero_n_2),
        .calc_bucket_set_addr_i_dld(calc_bucket_set_addr_i_dld),
        .calc_is_dummy_dld(calc_is_dummy_dld),
        .calc_is_zero_dld(calc_is_zero_dld),
        .clk(clk),
        .douta(mark_check_bucket_flag_out),
        .\gen_rd_a.gen_douta_pipe.gen_stages.douta_pipe_reg[1][0] (i_shiftreg_calc_bucket_set_addr_n_3),
        .processing_first_accept_flag(processing_first_accept_flag),
        .prsi_index_i(prsi_index_i));
  ponos_shiftreg_0 i_shiftreg_calc_is_dummy
       (.calc_is_dummy_dld(calc_is_dummy_dld),
        .clk(clk),
        .prsi_index_i(prsi_index_i));
  ponos_shiftreg_1 i_shiftreg_calc_is_zero
       (.\DELAY_BLOCK[3].shift_array_reg[4][0]_0 (i_shiftreg_calc_is_zero_n_1),
        .\DELAY_BLOCK[3].shift_array_reg[4][0]_1 (i_shiftreg_calc_is_zero_n_2),
        .\DELAY_BLOCK[3].shift_array_reg[4][0]_2 (i_shiftreg_calc_is_zero_n_3),
        .\DELAY_BLOCK[3].shift_array_reg[4][0]_3 (i_shiftreg_calc_is_zero_n_4),
        .\DELAY_BLOCK[3].shift_array_reg[4][0]_4 (i_shiftreg_calc_is_zero_n_5),
        .Q(\valid_dld_reg_n_0_[3] ),
        .acc_valid_o0(acc_valid_o0),
        .accept_flags_o({accept_flags_o[6],accept_flags_o[4:3],accept_flags_o[1]}),
        .\accept_flags_o_reg[1] (i_shiftreg_calc_bucket_set_addr_n_9),
        .\accept_flags_o_reg[3] (i_shiftreg_calc_bucket_set_addr_n_8),
        .\accept_flags_o_reg[4] (i_shiftreg_calc_bucket_set_addr_n_7),
        .\accept_flags_o_reg[6] (i_shiftreg_calc_bucket_set_addr_n_6),
        .calc_is_dummy_dld(calc_is_dummy_dld),
        .calc_is_zero(calc_is_zero),
        .calc_is_zero_dld(calc_is_zero_dld),
        .clk(clk),
        .douta(mark_check_bucket_flag_out),
        .processing_first_accept_flag(processing_first_accept_flag));
  ponos_shiftreg__parameterized2 i_shiftreg_point
       (.acc_point_o(acc_point_o),
        .clk(clk),
        .prsi_point_i(prsi_point_i));
  (* ADDR_WIDTH_A = "15" *) 
  (* ADDR_WIDTH_B = "15" *) 
  (* AUTO_SLEEP_TIME = "0" *) 
  (* BYTE_WRITE_WIDTH_A = "1" *) 
  (* BYTE_WRITE_WIDTH_B = "1" *) 
  (* CASCADE_HEIGHT = "0" *) 
  (* CLOCKING_MODE = "0" *) 
  (* ECC_BIT_RANGE = "[7:0]" *) 
  (* ECC_MODE = "0" *) 
  (* ECC_TYPE = "NONE" *) 
  (* IGNORE_INIT_SYNTH = "0" *) 
  (* MEMORY_INIT_FILE = "none" *) 
  (* MEMORY_INIT_PARAM = "" *) 
  (* MEMORY_OPTIMIZATION = "true" *) 
  (* MEMORY_PRIMITIVE = "0" *) 
  (* MEMORY_SIZE = "32768" *) 
  (* MESSAGE_CONTROL = "0" *) 
  (* P_CLOCKING_MODE = "0" *) 
  (* P_ECC_MODE = "0" *) 
  (* P_MEMORY_OPTIMIZATION = "1" *) 
  (* P_MEMORY_PRIMITIVE = "2" *) 
  (* P_WAKEUP_TIME = "0" *) 
  (* P_WRITE_MODE_A = "1" *) 
  (* P_WRITE_MODE_B = "1" *) 
  (* RAM_DECOMP = "auto" *) 
  (* READ_DATA_WIDTH_A = "1" *) 
  (* READ_DATA_WIDTH_B = "1" *) 
  (* READ_LATENCY_A = "3" *) 
  (* READ_LATENCY_B = "3" *) 
  (* READ_RESET_VALUE_A = "0" *) 
  (* READ_RESET_VALUE_B = "0" *) 
  (* RST_MODE_A = "SYNC" *) 
  (* RST_MODE_B = "SYNC" *) 
  (* SIM_ASSERT_CHK = "0" *) 
  (* USE_EMBEDDED_CONSTRAINT = "0" *) 
  (* USE_MEM_INIT = "1" *) 
  (* USE_MEM_INIT_MMI = "0" *) 
  (* WAKEUP_TIME = "0" *) 
  (* WRITE_DATA_WIDTH_A = "1" *) 
  (* WRITE_DATA_WIDTH_B = "1" *) 
  (* WRITE_MODE_A = "read_first" *) 
  (* WRITE_MODE_B = "read_first" *) 
  (* WRITE_PROTECT = "1" *) 
  (* XPM_MODULE = "TRUE" *) 
  ponos_xpm_memory_tdpram i_tdpram_flag_mem
       (.addra(mark_check_bucket_flag_addr),
        .addrb(clear_bucket_flag_addr),
        .clka(clk),
        .clkb(\<const0> ),
        .dina(\valid_dld_reg_n_0_[0] ),
        .dinb(\<const0> ),
        .douta(mark_check_bucket_flag_out),
        .ena(\<const1> ),
        .enb(\<const1> ),
        .injectdbiterra(\<const0> ),
        .injectdbiterrb(\<const0> ),
        .injectsbiterra(\<const0> ),
        .injectsbiterrb(\<const0> ),
        .regcea(\<const1> ),
        .regceb(\<const1> ),
        .rsta(prsi_ready_o_i_1_n_0),
        .rstb(\<const0> ),
        .sleep(\<const0> ),
        .wea(mark_check_bucket_flag_we),
        .web(clear_bucket_flag_we));
  FDRE #(
    .INIT(1'b0)) 
    \last_dld_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(prsi_last_i),
        .Q(\last_dld_reg_n_0_[0] ),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \last_dld_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\last_dld_reg_n_0_[0] ),
        .Q(\last_dld_reg_n_0_[1] ),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \last_dld_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\last_dld_reg_n_0_[1] ),
        .Q(\last_dld_reg_n_0_[2] ),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \last_dld_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\last_dld_reg_n_0_[2] ),
        .Q(\last_dld_reg_n_0_[3] ),
        .R(prsi_ready_o_i_1_n_0));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \mark_check_bucket_flag_addr[11]_i_1 
       (.I0(rst_n),
        .I1(prsi_ready_o),
        .I2(prsi_valid_i),
        .I3(i_shiftreg_calc_bucket_addr_n_13),
        .O(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \mark_check_bucket_flag_addr[12]_i_1 
       (.I0(prsi_valid_i),
        .I1(prsi_ready_o),
        .I2(rst_n),
        .I3(prsi_index_i[0]),
        .O(\mark_check_bucket_flag_addr[12]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \mark_check_bucket_flag_addr[13]_i_1 
       (.I0(prsi_valid_i),
        .I1(prsi_ready_o),
        .I2(rst_n),
        .I3(prsi_index_i[1]),
        .O(\mark_check_bucket_flag_addr[13]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \mark_check_bucket_flag_addr[14]_i_1 
       (.I0(prsi_valid_i),
        .I1(prsi_ready_o),
        .I2(rst_n),
        .I3(prsi_index_i[2]),
        .O(\mark_check_bucket_flag_addr[14]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[0]),
        .Q(mark_check_bucket_flag_addr[0]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[10]),
        .Q(mark_check_bucket_flag_addr[10]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[11]),
        .Q(mark_check_bucket_flag_addr[11]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\mark_check_bucket_flag_addr[12]_i_1_n_0 ),
        .Q(mark_check_bucket_flag_addr[12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\mark_check_bucket_flag_addr[13]_i_1_n_0 ),
        .Q(mark_check_bucket_flag_addr[13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\mark_check_bucket_flag_addr[14]_i_1_n_0 ),
        .Q(mark_check_bucket_flag_addr[14]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[1]),
        .Q(mark_check_bucket_flag_addr[1]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[2]),
        .Q(mark_check_bucket_flag_addr[2]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[3]),
        .Q(mark_check_bucket_flag_addr[3]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[4]),
        .Q(mark_check_bucket_flag_addr[4]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[5]),
        .Q(mark_check_bucket_flag_addr[5]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[6]),
        .Q(mark_check_bucket_flag_addr[6]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[7]),
        .Q(mark_check_bucket_flag_addr[7]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[8]),
        .Q(mark_check_bucket_flag_addr[8]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \mark_check_bucket_flag_addr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(data0[9]),
        .Q(mark_check_bucket_flag_addr[9]),
        .R(\mark_check_bucket_flag_addr[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hE0A00000)) 
    mark_check_bucket_flag_we_i_1
       (.I0(mark_check_bucket_flag_we_i_2_n_0),
        .I1(mark_check_bucket_flag_we_i_3_n_0),
        .I2(i_shiftreg_calc_bucket_addr_n_13),
        .I3(mark_check_bucket_flag_we_i_4_n_0),
        .I4(mark_check_bucket_flag_we_i_5_n_0),
        .O(mark_check_bucket_flag_we_i_1_n_0));
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'h6FF6)) 
    mark_check_bucket_flag_we_i_10
       (.I0(data0[1]),
        .I1(bm_bucket_addr_i[1]),
        .I2(data0[2]),
        .I3(bm_bucket_addr_i[2]),
        .O(mark_check_bucket_flag_we_i_10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT5 #(
    .INIT(32'h7DFFFF7D)) 
    mark_check_bucket_flag_we_i_11
       (.I0(bm_valid_i),
        .I1(bm_bucket_addr_i[11]),
        .I2(data0[11]),
        .I3(data0[0]),
        .I4(bm_bucket_addr_i[0]),
        .O(mark_check_bucket_flag_we_i_11_n_0));
  LUT6 #(
    .INIT(64'h31FF337DBEFFFFBE)) 
    mark_check_bucket_flag_we_i_2
       (.I0(bm_bucket_set_addr_i[0]),
        .I1(prsi_index_i[1]),
        .I2(bm_bucket_set_addr_i[1]),
        .I3(prsi_index_i[2]),
        .I4(bm_bucket_set_addr_i[2]),
        .I5(prsi_index_i[0]),
        .O(mark_check_bucket_flag_we_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    mark_check_bucket_flag_we_i_3
       (.I0(mark_check_bucket_flag_we_i_6_n_0),
        .I1(mark_check_bucket_flag_we_i_7_n_0),
        .I2(mark_check_bucket_flag_we_i_8_n_0),
        .I3(mark_check_bucket_flag_we_i_9_n_0),
        .I4(mark_check_bucket_flag_we_i_10_n_0),
        .I5(mark_check_bucket_flag_we_i_11_n_0),
        .O(mark_check_bucket_flag_we_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    mark_check_bucket_flag_we_i_4
       (.I0(prsi_index_i[2]),
        .I1(prsi_index_i[1]),
        .I2(prsi_index_i[0]),
        .O(mark_check_bucket_flag_we_i_4_n_0));
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT3 #(
    .INIT(8'h80)) 
    mark_check_bucket_flag_we_i_5
       (.I0(rst_n),
        .I1(prsi_ready_o),
        .I2(prsi_valid_i),
        .O(mark_check_bucket_flag_we_i_5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'h6FF6)) 
    mark_check_bucket_flag_we_i_6
       (.I0(data0[7]),
        .I1(bm_bucket_addr_i[7]),
        .I2(data0[8]),
        .I3(bm_bucket_addr_i[8]),
        .O(mark_check_bucket_flag_we_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT4 #(
    .INIT(16'h6FF6)) 
    mark_check_bucket_flag_we_i_7
       (.I0(data0[9]),
        .I1(bm_bucket_addr_i[9]),
        .I2(data0[10]),
        .I3(bm_bucket_addr_i[10]),
        .O(mark_check_bucket_flag_we_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT4 #(
    .INIT(16'h6FF6)) 
    mark_check_bucket_flag_we_i_8
       (.I0(data0[3]),
        .I1(bm_bucket_addr_i[3]),
        .I2(data0[4]),
        .I3(bm_bucket_addr_i[4]),
        .O(mark_check_bucket_flag_we_i_8_n_0));
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'h6FF6)) 
    mark_check_bucket_flag_we_i_9
       (.I0(data0[5]),
        .I1(bm_bucket_addr_i[5]),
        .I2(data0[6]),
        .I3(bm_bucket_addr_i[6]),
        .O(mark_check_bucket_flag_we_i_9_n_0));
  FDRE #(
    .INIT(1'b0)) 
    mark_check_bucket_flag_we_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(mark_check_bucket_flag_we_i_1_n_0),
        .Q(mark_check_bucket_flag_we),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hB8)) 
    processing_first_accept_flag_i_1
       (.I0(\last_dld_reg_n_0_[3] ),
        .I1(\valid_dld_reg_n_0_[3] ),
        .I2(processing_first_accept_flag),
        .O(processing_first_accept_flag_i_1_n_0));
  FDSE #(
    .INIT(1'b1)) 
    processing_first_accept_flag_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(processing_first_accept_flag_i_1_n_0),
        .Q(processing_first_accept_flag),
        .S(prsi_ready_o_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    prsi_ready_o_i_1
       (.I0(rst_n),
        .O(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    prsi_ready_o_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(init_done_i),
        .Q(prsi_ready_o),
        .R(prsi_ready_o_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    \valid_dld[0]_i_1 
       (.I0(prsi_ready_o),
        .I1(prsi_valid_i),
        .O(p_7_in));
  FDRE #(
    .INIT(1'b0)) 
    \valid_dld_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_7_in),
        .Q(\valid_dld_reg_n_0_[0] ),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \valid_dld_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\valid_dld_reg_n_0_[0] ),
        .Q(\valid_dld_reg_n_0_[1] ),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \valid_dld_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\valid_dld_reg_n_0_[1] ),
        .Q(\valid_dld_reg_n_0_[2] ),
        .R(prsi_ready_o_i_1_n_0));
  FDRE #(
    .INIT(1'b0)) 
    \valid_dld_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\valid_dld_reg_n_0_[2] ),
        .Q(\valid_dld_reg_n_0_[3] ),
        .R(prsi_ready_o_i_1_n_0));
endmodule
